LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;
USE IEEE.NUMERIC_STD.all;

ENTITY ENCODER_READING IS
	GENERIC (width:POSITIVE:=16);
	PORT (CHANNEL_A_RIGHT_1 	: IN std_logic; 
			CHANNEL_A_RIGHT_2 	: IN std_logic;
			CHANNEL_A_LEFT_1 		: IN std_logic;
			CHANNEL_A_LEFT_2 		: IN std_logic;
			CHANNEL_B_RIGHT_1 	: IN std_logic; 
			CHANNEL_B_RIGHT_2 	: IN std_logic;
			CHANNEL_B_LEFT_1 		: IN std_logic;
			CHANNEL_B_LEFT_2 		: IN std_logic; 
         reset 					: IN std_logic; 
         enable					: IN std_logic; 
         LEFT_COUNT		 		: OUT std_logic_vector(width-1 DOWNTO 0);
			RIGHT_COUNT		 		: OUT std_logic_vector(width-1 DOWNTO 0)
	);
END ENCODER_READING;

ARCHITECTURE MAIN OF ENCODER_READING IS
	SIGNAL LEFT_TICKS_1  : SIGNED(width-1 DOWNTO 0) := (others => '0');
	SIGNAL LEFT_TICKS_2  : SIGNED(width-1 DOWNTO 0) := (others => '0');
	SIGNAL RIGHT_TICKS_1 : SIGNED(width-1 DOWNTO 0) := (others => '0');
	SIGNAL RIGHT_TICKS_2 : SIGNED(width-1 DOWNTO 0) := (others => '0');
	
	SIGNAL LEFT_XOR_1  	: STD_LOGIC := '0';
	SIGNAL RIGHT_XOR_1 	: STD_LOGIC := '0';
	SIGNAL LEFT_XOR_2  	: STD_LOGIC := '0';
	SIGNAL RIGHT_XOR_2 	: STD_LOGIC := '0';
	
BEGIN

	-- SEE https://cdn.sparkfun.com/datasheets/Robotics/How%20to%20use%20a%20quadrature%20encoder.pdf
	RIGHT_XOR_1 <= CHANNEL_A_RIGHT_1 XOR CHANNEL_B_RIGHT_1;
	RIGHT_XOR_2 <= CHANNEL_A_RIGHT_2 XOR CHANNEL_B_RIGHT_2;
	LEFT_XOR_1  <= CHANNEL_A_LEFT_1 	XOR CHANNEL_B_LEFT_1;
	LEFT_XOR_2  <= CHANNEL_A_LEFT_2 	XOR CHANNEL_B_LEFT_2;
	
	COUNT_TICKS_RIGHT_1 : PROCESS (CHANNEL_A_RIGHT_1, CHANNEL_B_RIGHT_1, reset) IS
	BEGIN
		IF reset = '1' THEN
			RIGHT_TICKS_1 <= (others => '0');
		ELSIF RISING_EDGE(CHANNEL_A_RIGHT_1) THEN
			IF enable='1' THEN
				RIGHT_TICKS_1 <= RIGHT_TICKS_1 + 1;
			END IF;
		END IF;
	END PROCESS;
	
	COUNT_TICKS_RIGHT_2 : PROCESS (CHANNEL_A_RIGHT_2, CHANNEL_B_RIGHT_2, reset) IS
	BEGIN
		IF reset = '1' THEN
			RIGHT_TICKS_2 <= (others => '0');
		ELSIF RISING_EDGE(CHANNEL_A_RIGHT_2) THEN
			IF enable='1' THEN
				RIGHT_TICKS_2 <= RIGHT_TICKS_2 + 1;
			END IF;
		END IF;
	END PROCESS;
	
	RIGHT_COUNT <= std_logic_vector((RIGHT_TICKS_1 + RIGHT_TICKS_2)/2);
	
	COUNT_TICKS_LEFT_1 : PROCESS (CHANNEL_A_LEFT_1, CHANNEL_B_LEFT_1, reset) IS
	BEGIN
		IF reset = '1' THEN
			LEFT_TICKS_1<= (others => '0');
		ELSIF RISING_EDGE(CHANNEL_A_LEFT_1) THEN
			IF enable='1' THEN
				LEFT_TICKS_1 <= LEFT_TICKS_1 + 1;
			END IF;
		END IF;
	END PROCESS;
	
	COUNT_TICKS_LEFT_2 : PROCESS (CHANNEL_A_LEFT_2, CHANNEL_B_LEFT_2, reset) IS
	BEGIN
		IF reset = '1' THEN
			LEFT_TICKS_2 <= (others => '0');
		ELSIF RISING_EDGE(CHANNEL_A_LEFT_1) THEN
			IF enable='1' THEN
				LEFT_TICKS_2 <= LEFT_TICKS_2 + 1;
			END IF;
		END IF;
	END PROCESS;
	
	LEFT_COUNT <= std_logic_vector((LEFT_TICKS_1 + LEFT_TICKS_2)/2);
	
END MAIN;