-- NIOS.vhd

-- Generated using ACDS version 13.1 162 at 2015.08.31.20:25:04

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity NIOS is
	port (
		clk_clk                        : in    std_logic                     := '0';             --              clk.clk
		reset_reset_n                  : in    std_logic                     := '0';             --            reset.reset_n
		sdram_addr                     : out   std_logic_vector(12 downto 0);                    --            sdram.addr
		sdram_ba                       : out   std_logic_vector(1 downto 0);                     --                 .ba
		sdram_cas_n                    : out   std_logic;                                        --                 .cas_n
		sdram_cke                      : out   std_logic;                                        --                 .cke
		sdram_cs_n                     : out   std_logic;                                        --                 .cs_n
		sdram_dq                       : inout std_logic_vector(15 downto 0) := (others => '0'); --                 .dq
		sdram_dqm                      : out   std_logic_vector(1 downto 0);                     --                 .dqm
		sdram_ras_n                    : out   std_logic;                                        --                 .ras_n
		sdram_we_n                     : out   std_logic;                                        --                 .we_n
		epcs_dclk                      : out   std_logic;                                        --             epcs.dclk
		epcs_sce                       : out   std_logic;                                        --                 .sce
		epcs_sdo                       : out   std_logic;                                        --                 .sdo
		epcs_data0                     : in    std_logic                     := '0';             --                 .data0
		led_export                     : out   std_logic_vector(7 downto 0);                     --              led.export
		sw_export                      : in    std_logic_vector(3 downto 0)  := (others => '0'); --               sw.export
		key_export                     : in    std_logic_vector(1 downto 0)  := (others => '0'); --              key.export
		acelerometro_spi_I2C_SDAT      : inout std_logic                     := '0';             -- acelerometro_spi.I2C_SDAT
		acelerometro_spi_I2C_SCLK      : out   std_logic;                                        --                 .I2C_SCLK
		acelerometro_spi_G_SENSOR_CS_N : out   std_logic;                                        --                 .G_SENSOR_CS_N
		acelerometro_spi_G_SENSOR_INT  : in    std_logic                     := '0';             --                 .G_SENSOR_INT
		adc_sclk                       : out   std_logic;                                        --              adc.sclk
		adc_cs_n                       : out   std_logic;                                        --                 .cs_n
		adc_dout                       : in    std_logic                     := '0';             --                 .dout
		adc_din                        : out   std_logic;                                        --                 .din
		encoder_int_export             : in    std_logic_vector(3 downto 0)  := (others => '0'); --      encoder_int.export
		encoder_normal_export          : in    std_logic_vector(3 downto 0)  := (others => '0'); --   encoder_normal.export
		motores_export                 : out   std_logic_vector(5 downto 0);                     --          motores.export
		pwm1_export                    : out   std_logic_vector(7 downto 0);                     --             pwm1.export
		pwm2_export                    : out   std_logic_vector(7 downto 0);                     --             pwm2.export
		ctrl_i2c_export                : out   std_logic_vector(6 downto 0);                     --         ctrl_i2c.export
		data_out_i2c_export            : out   std_logic_vector(7 downto 0);                     --     data_out_i2c.export
		data_in_i2c_export             : in    std_logic_vector(7 downto 0)  := (others => '0'); --      data_in_i2c.export
		flag_i2c_export                : in    std_logic_vector(1 downto 0)  := (others => '0'); --         flag_i2c.export
		gps_rxd                        : in    std_logic                     := '0';             --              gps.rxd
		gps_txd                        : out   std_logic;                                        --                 .txd
		xbee_rxd                       : in    std_logic                     := '0';             --             xbee.rxd
		xbee_txd                       : out   std_logic;                                        --                 .txd
		dist1_rxd                      : in    std_logic                     := '0';             --            dist1.rxd
		dist1_txd                      : out   std_logic;                                        --                 .txd
		dist2_rxd                      : in    std_logic                     := '0';             --            dist2.rxd
		dist2_txd                      : out   std_logic;                                        --                 .txd
		dist3_rxd                      : in    std_logic                     := '0';             --            dist3.rxd
		dist3_txd                      : out   std_logic;                                        --                 .txd
		dist4_rxd                      : in    std_logic                     := '0';             --            dist4.rxd
		dist4_txd                      : out   std_logic                                         --                 .txd
	);
end entity NIOS;

architecture rtl of NIOS is
	component NIOS_CPU is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(26 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(26 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			i_readdatavalid                       : in  std_logic                     := 'X';             -- readdatavalid
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component NIOS_CPU;

	component NIOS_sys_id is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component NIOS_sys_id;

	component NIOS_SDRAM is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(23 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component NIOS_SDRAM;

	component NIOS_EPCS is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			reset_req     : in  std_logic                     := 'X';             -- reset_req
			address       : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			dataavailable : out std_logic;                                        -- dataavailable
			endofpacket   : out std_logic;                                        -- endofpacket
			read_n        : in  std_logic                     := 'X';             -- read_n
			readdata      : out std_logic_vector(31 downto 0);                    -- readdata
			readyfordata  : out std_logic;                                        -- readyfordata
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			irq           : out std_logic;                                        -- irq
			dclk          : out std_logic;                                        -- export
			sce           : out std_logic;                                        -- export
			sdo           : out std_logic;                                        -- export
			data0         : in  std_logic                     := 'X'              -- export
		);
	end component NIOS_EPCS;

	component NIOS_sys_timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component NIOS_sys_timer;

	component NIOS_LED is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component NIOS_LED;

	component NIOS_SW is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(3 downto 0)  := (others => 'X')  -- export
		);
	end component NIOS_SW;

	component NIOS_KEY is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOS_KEY;

	component NIOS_JTAG is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component NIOS_JTAG;

	component NIOS_sys_pll is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			c1        : out std_logic;                                        -- clk
			areset    : in  std_logic                     := 'X';             -- export
			locked    : out std_logic;                                        -- export
			phasedone : out std_logic                                         -- export
		);
	end component NIOS_sys_pll;

	component NIOS_ACELEROMETRO_SPI is
		port (
			clk           : in    std_logic                    := 'X';             -- clk
			reset         : in    std_logic                    := 'X';             -- reset
			address       : in    std_logic                    := 'X';             -- address
			byteenable    : in    std_logic                    := 'X';             -- byteenable
			read          : in    std_logic                    := 'X';             -- read
			write         : in    std_logic                    := 'X';             -- write
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			waitrequest   : out   std_logic;                                       -- waitrequest
			irq           : out   std_logic;                                       -- irq
			I2C_SDAT      : inout std_logic                    := 'X';             -- export
			I2C_SCLK      : out   std_logic;                                       -- export
			G_SENSOR_CS_N : out   std_logic;                                       -- export
			G_SENSOR_INT  : in    std_logic                    := 'X'              -- export
		);
	end component NIOS_ACELEROMETRO_SPI;

	component NIOS_ADC_DE0 is
		port (
			clock       : in  std_logic                     := 'X';             -- clk
			reset       : in  std_logic                     := 'X';             -- reset
			write       : in  std_logic                     := 'X';             -- write
			readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			address     : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			waitrequest : out std_logic;                                        -- waitrequest
			read        : in  std_logic                     := 'X';             -- read
			adc_sclk    : out std_logic;                                        -- export
			adc_cs_n    : out std_logic;                                        -- export
			adc_dout    : in  std_logic                     := 'X';             -- export
			adc_din     : out std_logic                                         -- export
		);
	end component NIOS_ADC_DE0;

	component NIOS_ENCODER_INT is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component NIOS_ENCODER_INT;

	component NIOS_MOTORES is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(5 downto 0)                      -- export
		);
	end component NIOS_MOTORES;

	component NIOS_CTRL_I2C is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component NIOS_CTRL_I2C;

	component NIOS_DATA_IN_I2C is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component NIOS_DATA_IN_I2C;

	component NIOS_FLAG_I2C is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component NIOS_FLAG_I2C;

	component NIOS_GPS is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			address       : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			begintransfer : in  std_logic                     := 'X';             -- begintransfer
			chipselect    : in  std_logic                     := 'X';             -- chipselect
			read_n        : in  std_logic                     := 'X';             -- read_n
			write_n       : in  std_logic                     := 'X';             -- write_n
			writedata     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata      : out std_logic_vector(15 downto 0);                    -- readdata
			dataavailable : out std_logic;                                        -- dataavailable
			readyfordata  : out std_logic;                                        -- readyfordata
			rxd           : in  std_logic                     := 'X';             -- export
			txd           : out std_logic;                                        -- export
			irq           : out std_logic                                         -- irq
		);
	end component NIOS_GPS;

	component NIOS_mm_interconnect_0 is
		port (
			clk_50_clk_clk                                                   : in  std_logic                     := 'X';             -- clk
			ram_clk_clk_clk                                                  : in  std_logic                     := 'X';             -- clk
			sys_clk_clk_clk                                                  : in  std_logic                     := 'X';             -- clk
			CPU_reset_n_reset_bridge_in_reset_reset                          : in  std_logic                     := 'X';             -- reset
			EPCS_reset_reset_bridge_in_reset_reset                           : in  std_logic                     := 'X';             -- reset
			MOTORES_reset_reset_bridge_in_reset_reset                        : in  std_logic                     := 'X';             -- reset
			sys_pll_inclk_interface_reset_reset_bridge_in_reset_reset        : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                                          : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest                                      : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable                                       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                                             : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                                         : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_write                                            : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata                                        : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess                                      : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address                                   : in  std_logic_vector(26 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest                               : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read                                      : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata                                  : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_instruction_master_readdatavalid                             : out std_logic;                                        -- readdatavalid
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_write       : out std_logic;                                        -- write
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_read        : out std_logic;                                        -- read
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_readdata    : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_writedata   : out std_logic_vector(7 downto 0);                     -- writedata
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_byteenable  : out std_logic_vector(0 downto 0);                     -- byteenable
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			ADC_DE0_adc_slave_address                                        : out std_logic_vector(2 downto 0);                     -- address
			ADC_DE0_adc_slave_write                                          : out std_logic;                                        -- write
			ADC_DE0_adc_slave_read                                           : out std_logic;                                        -- read
			ADC_DE0_adc_slave_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ADC_DE0_adc_slave_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			ADC_DE0_adc_slave_waitrequest                                    : in  std_logic                     := 'X';             -- waitrequest
			CPU_jtag_debug_module_address                                    : out std_logic_vector(8 downto 0);                     -- address
			CPU_jtag_debug_module_write                                      : out std_logic;                                        -- write
			CPU_jtag_debug_module_read                                       : out std_logic;                                        -- read
			CPU_jtag_debug_module_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_jtag_debug_module_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_jtag_debug_module_byteenable                                 : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_jtag_debug_module_waitrequest                                : in  std_logic                     := 'X';             -- waitrequest
			CPU_jtag_debug_module_debugaccess                                : out std_logic;                                        -- debugaccess
			CTRL_I2C_s1_address                                              : out std_logic_vector(1 downto 0);                     -- address
			CTRL_I2C_s1_write                                                : out std_logic;                                        -- write
			CTRL_I2C_s1_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CTRL_I2C_s1_writedata                                            : out std_logic_vector(31 downto 0);                    -- writedata
			CTRL_I2C_s1_chipselect                                           : out std_logic;                                        -- chipselect
			DATA_IN_I2C_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			DATA_IN_I2C_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DATA_OUT_I2C_s1_address                                          : out std_logic_vector(1 downto 0);                     -- address
			DATA_OUT_I2C_s1_write                                            : out std_logic;                                        -- write
			DATA_OUT_I2C_s1_readdata                                         : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			DATA_OUT_I2C_s1_writedata                                        : out std_logic_vector(31 downto 0);                    -- writedata
			DATA_OUT_I2C_s1_chipselect                                       : out std_logic;                                        -- chipselect
			DIST1_s1_address                                                 : out std_logic_vector(2 downto 0);                     -- address
			DIST1_s1_write                                                   : out std_logic;                                        -- write
			DIST1_s1_read                                                    : out std_logic;                                        -- read
			DIST1_s1_readdata                                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			DIST1_s1_writedata                                               : out std_logic_vector(15 downto 0);                    -- writedata
			DIST1_s1_begintransfer                                           : out std_logic;                                        -- begintransfer
			DIST1_s1_chipselect                                              : out std_logic;                                        -- chipselect
			DIST2_s1_address                                                 : out std_logic_vector(2 downto 0);                     -- address
			DIST2_s1_write                                                   : out std_logic;                                        -- write
			DIST2_s1_read                                                    : out std_logic;                                        -- read
			DIST2_s1_readdata                                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			DIST2_s1_writedata                                               : out std_logic_vector(15 downto 0);                    -- writedata
			DIST2_s1_begintransfer                                           : out std_logic;                                        -- begintransfer
			DIST2_s1_chipselect                                              : out std_logic;                                        -- chipselect
			DIST3_s1_address                                                 : out std_logic_vector(2 downto 0);                     -- address
			DIST3_s1_write                                                   : out std_logic;                                        -- write
			DIST3_s1_read                                                    : out std_logic;                                        -- read
			DIST3_s1_readdata                                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			DIST3_s1_writedata                                               : out std_logic_vector(15 downto 0);                    -- writedata
			DIST3_s1_begintransfer                                           : out std_logic;                                        -- begintransfer
			DIST3_s1_chipselect                                              : out std_logic;                                        -- chipselect
			DIST4_s1_address                                                 : out std_logic_vector(2 downto 0);                     -- address
			DIST4_s1_write                                                   : out std_logic;                                        -- write
			DIST4_s1_read                                                    : out std_logic;                                        -- read
			DIST4_s1_readdata                                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			DIST4_s1_writedata                                               : out std_logic_vector(15 downto 0);                    -- writedata
			DIST4_s1_begintransfer                                           : out std_logic;                                        -- begintransfer
			DIST4_s1_chipselect                                              : out std_logic;                                        -- chipselect
			ENCODER_INT_s1_address                                           : out std_logic_vector(1 downto 0);                     -- address
			ENCODER_INT_s1_write                                             : out std_logic;                                        -- write
			ENCODER_INT_s1_readdata                                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			ENCODER_INT_s1_writedata                                         : out std_logic_vector(31 downto 0);                    -- writedata
			ENCODER_INT_s1_chipselect                                        : out std_logic;                                        -- chipselect
			ENCODER_NORMAL_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			ENCODER_NORMAL_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			EPCS_epcs_control_port_address                                   : out std_logic_vector(8 downto 0);                     -- address
			EPCS_epcs_control_port_write                                     : out std_logic;                                        -- write
			EPCS_epcs_control_port_read                                      : out std_logic;                                        -- read
			EPCS_epcs_control_port_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			EPCS_epcs_control_port_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			EPCS_epcs_control_port_chipselect                                : out std_logic;                                        -- chipselect
			FLAG_I2C_s1_address                                              : out std_logic_vector(1 downto 0);                     -- address
			FLAG_I2C_s1_readdata                                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			GPS_s1_address                                                   : out std_logic_vector(2 downto 0);                     -- address
			GPS_s1_write                                                     : out std_logic;                                        -- write
			GPS_s1_read                                                      : out std_logic;                                        -- read
			GPS_s1_readdata                                                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			GPS_s1_writedata                                                 : out std_logic_vector(15 downto 0);                    -- writedata
			GPS_s1_begintransfer                                             : out std_logic;                                        -- begintransfer
			GPS_s1_chipselect                                                : out std_logic;                                        -- chipselect
			JTAG_avalon_jtag_slave_address                                   : out std_logic_vector(0 downto 0);                     -- address
			JTAG_avalon_jtag_slave_write                                     : out std_logic;                                        -- write
			JTAG_avalon_jtag_slave_read                                      : out std_logic;                                        -- read
			JTAG_avalon_jtag_slave_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			JTAG_avalon_jtag_slave_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			JTAG_avalon_jtag_slave_waitrequest                               : in  std_logic                     := 'X';             -- waitrequest
			JTAG_avalon_jtag_slave_chipselect                                : out std_logic;                                        -- chipselect
			KEY_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			KEY_s1_write                                                     : out std_logic;                                        -- write
			KEY_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			KEY_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			KEY_s1_chipselect                                                : out std_logic;                                        -- chipselect
			LED_s1_address                                                   : out std_logic_vector(1 downto 0);                     -- address
			LED_s1_write                                                     : out std_logic;                                        -- write
			LED_s1_readdata                                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			LED_s1_writedata                                                 : out std_logic_vector(31 downto 0);                    -- writedata
			LED_s1_chipselect                                                : out std_logic;                                        -- chipselect
			MOTORES_s1_address                                               : out std_logic_vector(1 downto 0);                     -- address
			MOTORES_s1_write                                                 : out std_logic;                                        -- write
			MOTORES_s1_readdata                                              : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			MOTORES_s1_writedata                                             : out std_logic_vector(31 downto 0);                    -- writedata
			MOTORES_s1_chipselect                                            : out std_logic;                                        -- chipselect
			PWM1_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			PWM1_s1_write                                                    : out std_logic;                                        -- write
			PWM1_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PWM1_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			PWM1_s1_chipselect                                               : out std_logic;                                        -- chipselect
			PWM2_s1_address                                                  : out std_logic_vector(1 downto 0);                     -- address
			PWM2_s1_write                                                    : out std_logic;                                        -- write
			PWM2_s1_readdata                                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			PWM2_s1_writedata                                                : out std_logic_vector(31 downto 0);                    -- writedata
			PWM2_s1_chipselect                                               : out std_logic;                                        -- chipselect
			SDRAM_s1_address                                                 : out std_logic_vector(23 downto 0);                    -- address
			SDRAM_s1_write                                                   : out std_logic;                                        -- write
			SDRAM_s1_read                                                    : out std_logic;                                        -- read
			SDRAM_s1_readdata                                                : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SDRAM_s1_writedata                                               : out std_logic_vector(15 downto 0);                    -- writedata
			SDRAM_s1_byteenable                                              : out std_logic_vector(1 downto 0);                     -- byteenable
			SDRAM_s1_readdatavalid                                           : in  std_logic                     := 'X';             -- readdatavalid
			SDRAM_s1_waitrequest                                             : in  std_logic                     := 'X';             -- waitrequest
			SDRAM_s1_chipselect                                              : out std_logic;                                        -- chipselect
			SW_s1_address                                                    : out std_logic_vector(1 downto 0);                     -- address
			SW_s1_readdata                                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sys_id_control_slave_address                                     : out std_logic_vector(0 downto 0);                     -- address
			sys_id_control_slave_readdata                                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sys_pll_pll_slave_address                                        : out std_logic_vector(1 downto 0);                     -- address
			sys_pll_pll_slave_write                                          : out std_logic;                                        -- write
			sys_pll_pll_slave_read                                           : out std_logic;                                        -- read
			sys_pll_pll_slave_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sys_pll_pll_slave_writedata                                      : out std_logic_vector(31 downto 0);                    -- writedata
			sys_timer_s1_address                                             : out std_logic_vector(2 downto 0);                     -- address
			sys_timer_s1_write                                               : out std_logic;                                        -- write
			sys_timer_s1_readdata                                            : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sys_timer_s1_writedata                                           : out std_logic_vector(15 downto 0);                    -- writedata
			sys_timer_s1_chipselect                                          : out std_logic;                                        -- chipselect
			XBEE_s1_address                                                  : out std_logic_vector(2 downto 0);                     -- address
			XBEE_s1_write                                                    : out std_logic;                                        -- write
			XBEE_s1_read                                                     : out std_logic;                                        -- read
			XBEE_s1_readdata                                                 : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			XBEE_s1_writedata                                                : out std_logic_vector(15 downto 0);                    -- writedata
			XBEE_s1_begintransfer                                            : out std_logic;                                        -- begintransfer
			XBEE_s1_chipselect                                               : out std_logic                                         -- chipselect
		);
	end component NIOS_mm_interconnect_0;

	component NIOS_irq_mapper is
		port (
			clk            : in  std_logic                     := 'X'; -- clk
			reset          : in  std_logic                     := 'X'; -- reset
			receiver0_irq  : in  std_logic                     := 'X'; -- irq
			receiver1_irq  : in  std_logic                     := 'X'; -- irq
			receiver2_irq  : in  std_logic                     := 'X'; -- irq
			receiver3_irq  : in  std_logic                     := 'X'; -- irq
			receiver4_irq  : in  std_logic                     := 'X'; -- irq
			receiver5_irq  : in  std_logic                     := 'X'; -- irq
			receiver6_irq  : in  std_logic                     := 'X'; -- irq
			receiver7_irq  : in  std_logic                     := 'X'; -- irq
			receiver8_irq  : in  std_logic                     := 'X'; -- irq
			receiver9_irq  : in  std_logic                     := 'X'; -- irq
			receiver10_irq : in  std_logic                     := 'X'; -- irq
			receiver11_irq : in  std_logic                     := 'X'; -- irq
			sender_irq     : out std_logic_vector(31 downto 0)         -- irq
		);
	end component NIOS_irq_mapper;

	component nios_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_rst_controller;

	component nios_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_rst_controller_001;

	component nios_rst_controller_002 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_in1      : in  std_logic := 'X'; -- reset
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component nios_rst_controller_002;

	signal sys_pll_c0_clk                                                                     : std_logic;                     -- sys_pll:c0 -> [ACELEROMETRO_SPI:clk, ADC_DE0:clock, CPU:clk, CTRL_I2C:clk, DATA_IN_I2C:clk, DATA_OUT_I2C:clk, DIST1:clk, DIST2:clk, DIST3:clk, DIST4:clk, ENCODER_INT:clk, ENCODER_NORMAL:clk, EPCS:clk, FLAG_I2C:clk, GPS:clk, JTAG:clk, KEY:clk, LED:clk, PWM1:clk, PWM2:clk, SDRAM:clk, SW:clk, XBEE:clk, irq_mapper:clk, mm_interconnect_0:sys_clk_clk_clk, rst_controller:clk, rst_controller_001:clk, sys_id:clock, sys_timer:clk]
	signal sys_pll_c1_clk                                                                     : std_logic;                     -- sys_pll:c1 -> [MOTORES:clk, mm_interconnect_0:ram_clk_clk_clk, rst_controller_003:clk]
	signal mm_interconnect_0_led_s1_writedata                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:LED_s1_writedata -> LED:writedata
	signal mm_interconnect_0_led_s1_address                                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:LED_s1_address -> LED:address
	signal mm_interconnect_0_led_s1_chipselect                                                : std_logic;                     -- mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	signal mm_interconnect_0_led_s1_write                                                     : std_logic;                     -- mm_interconnect_0:LED_s1_write -> mm_interconnect_0_led_s1_write:in
	signal mm_interconnect_0_led_s1_readdata                                                  : std_logic_vector(31 downto 0); -- LED:readdata -> mm_interconnect_0:LED_s1_readdata
	signal mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_waitrequest : std_logic;                     -- ACELEROMETRO_SPI:waitrequest -> mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_waitrequest
	signal mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_writedata   : std_logic_vector(7 downto 0);  -- mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_writedata -> ACELEROMETRO_SPI:writedata
	signal mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_address     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_address -> ACELEROMETRO_SPI:address
	signal mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_write       : std_logic;                     -- mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_write -> ACELEROMETRO_SPI:write
	signal mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_read        : std_logic;                     -- mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_read -> ACELEROMETRO_SPI:read
	signal mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_readdata    : std_logic_vector(7 downto 0);  -- ACELEROMETRO_SPI:readdata -> mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_readdata
	signal mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_byteenable  : std_logic_vector(0 downto 0);  -- mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_byteenable -> ACELEROMETRO_SPI:byteenable
	signal mm_interconnect_0_pwm2_s1_writedata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:PWM2_s1_writedata -> PWM2:writedata
	signal mm_interconnect_0_pwm2_s1_address                                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PWM2_s1_address -> PWM2:address
	signal mm_interconnect_0_pwm2_s1_chipselect                                               : std_logic;                     -- mm_interconnect_0:PWM2_s1_chipselect -> PWM2:chipselect
	signal mm_interconnect_0_pwm2_s1_write                                                    : std_logic;                     -- mm_interconnect_0:PWM2_s1_write -> mm_interconnect_0_pwm2_s1_write:in
	signal mm_interconnect_0_pwm2_s1_readdata                                                 : std_logic_vector(31 downto 0); -- PWM2:readdata -> mm_interconnect_0:PWM2_s1_readdata
	signal mm_interconnect_0_dist1_s1_writedata                                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:DIST1_s1_writedata -> DIST1:writedata
	signal mm_interconnect_0_dist1_s1_address                                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:DIST1_s1_address -> DIST1:address
	signal mm_interconnect_0_dist1_s1_chipselect                                              : std_logic;                     -- mm_interconnect_0:DIST1_s1_chipselect -> DIST1:chipselect
	signal mm_interconnect_0_dist1_s1_write                                                   : std_logic;                     -- mm_interconnect_0:DIST1_s1_write -> mm_interconnect_0_dist1_s1_write:in
	signal mm_interconnect_0_dist1_s1_read                                                    : std_logic;                     -- mm_interconnect_0:DIST1_s1_read -> mm_interconnect_0_dist1_s1_read:in
	signal mm_interconnect_0_dist1_s1_readdata                                                : std_logic_vector(15 downto 0); -- DIST1:readdata -> mm_interconnect_0:DIST1_s1_readdata
	signal mm_interconnect_0_dist1_s1_begintransfer                                           : std_logic;                     -- mm_interconnect_0:DIST1_s1_begintransfer -> DIST1:begintransfer
	signal mm_interconnect_0_sys_id_control_slave_address                                     : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	signal mm_interconnect_0_sys_id_control_slave_readdata                                    : std_logic_vector(31 downto 0); -- sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	signal mm_interconnect_0_gps_s1_writedata                                                 : std_logic_vector(15 downto 0); -- mm_interconnect_0:GPS_s1_writedata -> GPS:writedata
	signal mm_interconnect_0_gps_s1_address                                                   : std_logic_vector(2 downto 0);  -- mm_interconnect_0:GPS_s1_address -> GPS:address
	signal mm_interconnect_0_gps_s1_chipselect                                                : std_logic;                     -- mm_interconnect_0:GPS_s1_chipselect -> GPS:chipselect
	signal mm_interconnect_0_gps_s1_write                                                     : std_logic;                     -- mm_interconnect_0:GPS_s1_write -> mm_interconnect_0_gps_s1_write:in
	signal mm_interconnect_0_gps_s1_read                                                      : std_logic;                     -- mm_interconnect_0:GPS_s1_read -> mm_interconnect_0_gps_s1_read:in
	signal mm_interconnect_0_gps_s1_readdata                                                  : std_logic_vector(15 downto 0); -- GPS:readdata -> mm_interconnect_0:GPS_s1_readdata
	signal mm_interconnect_0_gps_s1_begintransfer                                             : std_logic;                     -- mm_interconnect_0:GPS_s1_begintransfer -> GPS:begintransfer
	signal mm_interconnect_0_dist3_s1_writedata                                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:DIST3_s1_writedata -> DIST3:writedata
	signal mm_interconnect_0_dist3_s1_address                                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:DIST3_s1_address -> DIST3:address
	signal mm_interconnect_0_dist3_s1_chipselect                                              : std_logic;                     -- mm_interconnect_0:DIST3_s1_chipselect -> DIST3:chipselect
	signal mm_interconnect_0_dist3_s1_write                                                   : std_logic;                     -- mm_interconnect_0:DIST3_s1_write -> mm_interconnect_0_dist3_s1_write:in
	signal mm_interconnect_0_dist3_s1_read                                                    : std_logic;                     -- mm_interconnect_0:DIST3_s1_read -> mm_interconnect_0_dist3_s1_read:in
	signal mm_interconnect_0_dist3_s1_readdata                                                : std_logic_vector(15 downto 0); -- DIST3:readdata -> mm_interconnect_0:DIST3_s1_readdata
	signal mm_interconnect_0_dist3_s1_begintransfer                                           : std_logic;                     -- mm_interconnect_0:DIST3_s1_begintransfer -> DIST3:begintransfer
	signal mm_interconnect_0_epcs_epcs_control_port_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:EPCS_epcs_control_port_writedata -> EPCS:writedata
	signal mm_interconnect_0_epcs_epcs_control_port_address                                   : std_logic_vector(8 downto 0);  -- mm_interconnect_0:EPCS_epcs_control_port_address -> EPCS:address
	signal mm_interconnect_0_epcs_epcs_control_port_chipselect                                : std_logic;                     -- mm_interconnect_0:EPCS_epcs_control_port_chipselect -> EPCS:chipselect
	signal mm_interconnect_0_epcs_epcs_control_port_write                                     : std_logic;                     -- mm_interconnect_0:EPCS_epcs_control_port_write -> mm_interconnect_0_epcs_epcs_control_port_write:in
	signal mm_interconnect_0_epcs_epcs_control_port_read                                      : std_logic;                     -- mm_interconnect_0:EPCS_epcs_control_port_read -> mm_interconnect_0_epcs_epcs_control_port_read:in
	signal mm_interconnect_0_epcs_epcs_control_port_readdata                                  : std_logic_vector(31 downto 0); -- EPCS:readdata -> mm_interconnect_0:EPCS_epcs_control_port_readdata
	signal mm_interconnect_0_sw_s1_address                                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SW_s1_address -> SW:address
	signal mm_interconnect_0_sw_s1_readdata                                                   : std_logic_vector(31 downto 0); -- SW:readdata -> mm_interconnect_0:SW_s1_readdata
	signal mm_interconnect_0_xbee_s1_writedata                                                : std_logic_vector(15 downto 0); -- mm_interconnect_0:XBEE_s1_writedata -> XBEE:writedata
	signal mm_interconnect_0_xbee_s1_address                                                  : std_logic_vector(2 downto 0);  -- mm_interconnect_0:XBEE_s1_address -> XBEE:address
	signal mm_interconnect_0_xbee_s1_chipselect                                               : std_logic;                     -- mm_interconnect_0:XBEE_s1_chipselect -> XBEE:chipselect
	signal mm_interconnect_0_xbee_s1_write                                                    : std_logic;                     -- mm_interconnect_0:XBEE_s1_write -> mm_interconnect_0_xbee_s1_write:in
	signal mm_interconnect_0_xbee_s1_read                                                     : std_logic;                     -- mm_interconnect_0:XBEE_s1_read -> mm_interconnect_0_xbee_s1_read:in
	signal mm_interconnect_0_xbee_s1_readdata                                                 : std_logic_vector(15 downto 0); -- XBEE:readdata -> mm_interconnect_0:XBEE_s1_readdata
	signal mm_interconnect_0_xbee_s1_begintransfer                                            : std_logic;                     -- mm_interconnect_0:XBEE_s1_begintransfer -> XBEE:begintransfer
	signal mm_interconnect_0_sys_timer_s1_writedata                                           : std_logic_vector(15 downto 0); -- mm_interconnect_0:sys_timer_s1_writedata -> sys_timer:writedata
	signal mm_interconnect_0_sys_timer_s1_address                                             : std_logic_vector(2 downto 0);  -- mm_interconnect_0:sys_timer_s1_address -> sys_timer:address
	signal mm_interconnect_0_sys_timer_s1_chipselect                                          : std_logic;                     -- mm_interconnect_0:sys_timer_s1_chipselect -> sys_timer:chipselect
	signal mm_interconnect_0_sys_timer_s1_write                                               : std_logic;                     -- mm_interconnect_0:sys_timer_s1_write -> mm_interconnect_0_sys_timer_s1_write:in
	signal mm_interconnect_0_sys_timer_s1_readdata                                            : std_logic_vector(15 downto 0); -- sys_timer:readdata -> mm_interconnect_0:sys_timer_s1_readdata
	signal mm_interconnect_0_encoder_int_s1_writedata                                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:ENCODER_INT_s1_writedata -> ENCODER_INT:writedata
	signal mm_interconnect_0_encoder_int_s1_address                                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ENCODER_INT_s1_address -> ENCODER_INT:address
	signal mm_interconnect_0_encoder_int_s1_chipselect                                        : std_logic;                     -- mm_interconnect_0:ENCODER_INT_s1_chipselect -> ENCODER_INT:chipselect
	signal mm_interconnect_0_encoder_int_s1_write                                             : std_logic;                     -- mm_interconnect_0:ENCODER_INT_s1_write -> mm_interconnect_0_encoder_int_s1_write:in
	signal mm_interconnect_0_encoder_int_s1_readdata                                          : std_logic_vector(31 downto 0); -- ENCODER_INT:readdata -> mm_interconnect_0:ENCODER_INT_s1_readdata
	signal mm_interconnect_0_dist4_s1_writedata                                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:DIST4_s1_writedata -> DIST4:writedata
	signal mm_interconnect_0_dist4_s1_address                                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:DIST4_s1_address -> DIST4:address
	signal mm_interconnect_0_dist4_s1_chipselect                                              : std_logic;                     -- mm_interconnect_0:DIST4_s1_chipselect -> DIST4:chipselect
	signal mm_interconnect_0_dist4_s1_write                                                   : std_logic;                     -- mm_interconnect_0:DIST4_s1_write -> mm_interconnect_0_dist4_s1_write:in
	signal mm_interconnect_0_dist4_s1_read                                                    : std_logic;                     -- mm_interconnect_0:DIST4_s1_read -> mm_interconnect_0_dist4_s1_read:in
	signal mm_interconnect_0_dist4_s1_readdata                                                : std_logic_vector(15 downto 0); -- DIST4:readdata -> mm_interconnect_0:DIST4_s1_readdata
	signal mm_interconnect_0_dist4_s1_begintransfer                                           : std_logic;                     -- mm_interconnect_0:DIST4_s1_begintransfer -> DIST4:begintransfer
	signal mm_interconnect_0_cpu_jtag_debug_module_waitrequest                                : std_logic;                     -- CPU:jtag_debug_module_waitrequest -> mm_interconnect_0:CPU_jtag_debug_module_waitrequest
	signal mm_interconnect_0_cpu_jtag_debug_module_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	signal mm_interconnect_0_cpu_jtag_debug_module_address                                    : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	signal mm_interconnect_0_cpu_jtag_debug_module_write                                      : std_logic;                     -- mm_interconnect_0:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	signal mm_interconnect_0_cpu_jtag_debug_module_read                                       : std_logic;                     -- mm_interconnect_0:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	signal mm_interconnect_0_cpu_jtag_debug_module_readdata                                   : std_logic_vector(31 downto 0); -- CPU:jtag_debug_module_readdata -> mm_interconnect_0:CPU_jtag_debug_module_readdata
	signal mm_interconnect_0_cpu_jtag_debug_module_debugaccess                                : std_logic;                     -- mm_interconnect_0:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	signal mm_interconnect_0_cpu_jtag_debug_module_byteenable                                 : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	signal mm_interconnect_0_data_out_i2c_s1_writedata                                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:DATA_OUT_I2C_s1_writedata -> DATA_OUT_I2C:writedata
	signal mm_interconnect_0_data_out_i2c_s1_address                                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:DATA_OUT_I2C_s1_address -> DATA_OUT_I2C:address
	signal mm_interconnect_0_data_out_i2c_s1_chipselect                                       : std_logic;                     -- mm_interconnect_0:DATA_OUT_I2C_s1_chipselect -> DATA_OUT_I2C:chipselect
	signal mm_interconnect_0_data_out_i2c_s1_write                                            : std_logic;                     -- mm_interconnect_0:DATA_OUT_I2C_s1_write -> mm_interconnect_0_data_out_i2c_s1_write:in
	signal mm_interconnect_0_data_out_i2c_s1_readdata                                         : std_logic_vector(31 downto 0); -- DATA_OUT_I2C:readdata -> mm_interconnect_0:DATA_OUT_I2C_s1_readdata
	signal mm_interconnect_0_key_s1_writedata                                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:KEY_s1_writedata -> KEY:writedata
	signal mm_interconnect_0_key_s1_address                                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:KEY_s1_address -> KEY:address
	signal mm_interconnect_0_key_s1_chipselect                                                : std_logic;                     -- mm_interconnect_0:KEY_s1_chipselect -> KEY:chipselect
	signal mm_interconnect_0_key_s1_write                                                     : std_logic;                     -- mm_interconnect_0:KEY_s1_write -> mm_interconnect_0_key_s1_write:in
	signal mm_interconnect_0_key_s1_readdata                                                  : std_logic_vector(31 downto 0); -- KEY:readdata -> mm_interconnect_0:KEY_s1_readdata
	signal mm_interconnect_0_data_in_i2c_s1_address                                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:DATA_IN_I2C_s1_address -> DATA_IN_I2C:address
	signal mm_interconnect_0_data_in_i2c_s1_readdata                                          : std_logic_vector(31 downto 0); -- DATA_IN_I2C:readdata -> mm_interconnect_0:DATA_IN_I2C_s1_readdata
	signal mm_interconnect_0_sys_pll_pll_slave_writedata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:sys_pll_pll_slave_writedata -> sys_pll:writedata
	signal mm_interconnect_0_sys_pll_pll_slave_address                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sys_pll_pll_slave_address -> sys_pll:address
	signal mm_interconnect_0_sys_pll_pll_slave_write                                          : std_logic;                     -- mm_interconnect_0:sys_pll_pll_slave_write -> sys_pll:write
	signal mm_interconnect_0_sys_pll_pll_slave_read                                           : std_logic;                     -- mm_interconnect_0:sys_pll_pll_slave_read -> sys_pll:read
	signal mm_interconnect_0_sys_pll_pll_slave_readdata                                       : std_logic_vector(31 downto 0); -- sys_pll:readdata -> mm_interconnect_0:sys_pll_pll_slave_readdata
	signal cpu_data_master_waitrequest                                                        : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_writedata                                                          : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_data_master_address                                                            : std_logic_vector(26 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_write                                                              : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_read                                                               : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_readdata                                                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_debugaccess                                                        : std_logic;                     -- CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_byteenable                                                         : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal mm_interconnect_0_ctrl_i2c_s1_writedata                                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:CTRL_I2C_s1_writedata -> CTRL_I2C:writedata
	signal mm_interconnect_0_ctrl_i2c_s1_address                                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:CTRL_I2C_s1_address -> CTRL_I2C:address
	signal mm_interconnect_0_ctrl_i2c_s1_chipselect                                           : std_logic;                     -- mm_interconnect_0:CTRL_I2C_s1_chipselect -> CTRL_I2C:chipselect
	signal mm_interconnect_0_ctrl_i2c_s1_write                                                : std_logic;                     -- mm_interconnect_0:CTRL_I2C_s1_write -> mm_interconnect_0_ctrl_i2c_s1_write:in
	signal mm_interconnect_0_ctrl_i2c_s1_readdata                                             : std_logic_vector(31 downto 0); -- CTRL_I2C:readdata -> mm_interconnect_0:CTRL_I2C_s1_readdata
	signal cpu_instruction_master_waitrequest                                                 : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                                     : std_logic_vector(26 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                                        : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal cpu_instruction_master_readdata                                                    : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_instruction_master_readdatavalid                                               : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	signal mm_interconnect_0_flag_i2c_s1_address                                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:FLAG_I2C_s1_address -> FLAG_I2C:address
	signal mm_interconnect_0_flag_i2c_s1_readdata                                             : std_logic_vector(31 downto 0); -- FLAG_I2C:readdata -> mm_interconnect_0:FLAG_I2C_s1_readdata
	signal mm_interconnect_0_encoder_normal_s1_address                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:ENCODER_NORMAL_s1_address -> ENCODER_NORMAL:address
	signal mm_interconnect_0_encoder_normal_s1_readdata                                       : std_logic_vector(31 downto 0); -- ENCODER_NORMAL:readdata -> mm_interconnect_0:ENCODER_NORMAL_s1_readdata
	signal mm_interconnect_0_motores_s1_writedata                                             : std_logic_vector(31 downto 0); -- mm_interconnect_0:MOTORES_s1_writedata -> MOTORES:writedata
	signal mm_interconnect_0_motores_s1_address                                               : std_logic_vector(1 downto 0);  -- mm_interconnect_0:MOTORES_s1_address -> MOTORES:address
	signal mm_interconnect_0_motores_s1_chipselect                                            : std_logic;                     -- mm_interconnect_0:MOTORES_s1_chipselect -> MOTORES:chipselect
	signal mm_interconnect_0_motores_s1_write                                                 : std_logic;                     -- mm_interconnect_0:MOTORES_s1_write -> mm_interconnect_0_motores_s1_write:in
	signal mm_interconnect_0_motores_s1_readdata                                              : std_logic_vector(31 downto 0); -- MOTORES:readdata -> mm_interconnect_0:MOTORES_s1_readdata
	signal mm_interconnect_0_adc_de0_adc_slave_waitrequest                                    : std_logic;                     -- ADC_DE0:waitrequest -> mm_interconnect_0:ADC_DE0_adc_slave_waitrequest
	signal mm_interconnect_0_adc_de0_adc_slave_writedata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:ADC_DE0_adc_slave_writedata -> ADC_DE0:writedata
	signal mm_interconnect_0_adc_de0_adc_slave_address                                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:ADC_DE0_adc_slave_address -> ADC_DE0:address
	signal mm_interconnect_0_adc_de0_adc_slave_write                                          : std_logic;                     -- mm_interconnect_0:ADC_DE0_adc_slave_write -> ADC_DE0:write
	signal mm_interconnect_0_adc_de0_adc_slave_read                                           : std_logic;                     -- mm_interconnect_0:ADC_DE0_adc_slave_read -> ADC_DE0:read
	signal mm_interconnect_0_adc_de0_adc_slave_readdata                                       : std_logic_vector(31 downto 0); -- ADC_DE0:readdata -> mm_interconnect_0:ADC_DE0_adc_slave_readdata
	signal mm_interconnect_0_pwm1_s1_writedata                                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:PWM1_s1_writedata -> PWM1:writedata
	signal mm_interconnect_0_pwm1_s1_address                                                  : std_logic_vector(1 downto 0);  -- mm_interconnect_0:PWM1_s1_address -> PWM1:address
	signal mm_interconnect_0_pwm1_s1_chipselect                                               : std_logic;                     -- mm_interconnect_0:PWM1_s1_chipselect -> PWM1:chipselect
	signal mm_interconnect_0_pwm1_s1_write                                                    : std_logic;                     -- mm_interconnect_0:PWM1_s1_write -> mm_interconnect_0_pwm1_s1_write:in
	signal mm_interconnect_0_pwm1_s1_readdata                                                 : std_logic_vector(31 downto 0); -- PWM1:readdata -> mm_interconnect_0:PWM1_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                             : std_logic;                     -- SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_writedata                                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	signal mm_interconnect_0_sdram_s1_address                                                 : std_logic_vector(23 downto 0); -- mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	signal mm_interconnect_0_sdram_s1_chipselect                                              : std_logic;                     -- mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	signal mm_interconnect_0_sdram_s1_write                                                   : std_logic;                     -- mm_interconnect_0:SDRAM_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_read                                                    : std_logic;                     -- mm_interconnect_0:SDRAM_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_readdata                                                : std_logic_vector(15 downto 0); -- SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	signal mm_interconnect_0_sdram_s1_readdatavalid                                           : std_logic;                     -- SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_byteenable                                              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SDRAM_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_dist2_s1_writedata                                               : std_logic_vector(15 downto 0); -- mm_interconnect_0:DIST2_s1_writedata -> DIST2:writedata
	signal mm_interconnect_0_dist2_s1_address                                                 : std_logic_vector(2 downto 0);  -- mm_interconnect_0:DIST2_s1_address -> DIST2:address
	signal mm_interconnect_0_dist2_s1_chipselect                                              : std_logic;                     -- mm_interconnect_0:DIST2_s1_chipselect -> DIST2:chipselect
	signal mm_interconnect_0_dist2_s1_write                                                   : std_logic;                     -- mm_interconnect_0:DIST2_s1_write -> mm_interconnect_0_dist2_s1_write:in
	signal mm_interconnect_0_dist2_s1_read                                                    : std_logic;                     -- mm_interconnect_0:DIST2_s1_read -> mm_interconnect_0_dist2_s1_read:in
	signal mm_interconnect_0_dist2_s1_readdata                                                : std_logic_vector(15 downto 0); -- DIST2:readdata -> mm_interconnect_0:DIST2_s1_readdata
	signal mm_interconnect_0_dist2_s1_begintransfer                                           : std_logic;                     -- mm_interconnect_0:DIST2_s1_begintransfer -> DIST2:begintransfer
	signal mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest                               : std_logic;                     -- JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_avalon_jtag_slave_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	signal mm_interconnect_0_jtag_avalon_jtag_slave_address                                   : std_logic_vector(0 downto 0);  -- mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	signal mm_interconnect_0_jtag_avalon_jtag_slave_chipselect                                : std_logic;                     -- mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write                                     : std_logic;                     -- mm_interconnect_0:JTAG_avalon_jtag_slave_write -> mm_interconnect_0_jtag_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read                                      : std_logic;                     -- mm_interconnect_0:JTAG_avalon_jtag_slave_read -> mm_interconnect_0_jtag_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_avalon_jtag_slave_readdata                                  : std_logic_vector(31 downto 0); -- JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	signal irq_mapper_receiver0_irq                                                           : std_logic;                     -- EPCS:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                           : std_logic;                     -- sys_timer:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                           : std_logic;                     -- JTAG:av_irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                                           : std_logic;                     -- KEY:irq -> irq_mapper:receiver3_irq
	signal irq_mapper_receiver4_irq                                                           : std_logic;                     -- ENCODER_INT:irq -> irq_mapper:receiver4_irq
	signal irq_mapper_receiver5_irq                                                           : std_logic;                     -- ACELEROMETRO_SPI:irq -> irq_mapper:receiver5_irq
	signal irq_mapper_receiver6_irq                                                           : std_logic;                     -- GPS:irq -> irq_mapper:receiver6_irq
	signal irq_mapper_receiver7_irq                                                           : std_logic;                     -- XBEE:irq -> irq_mapper:receiver7_irq
	signal irq_mapper_receiver8_irq                                                           : std_logic;                     -- DIST1:irq -> irq_mapper:receiver8_irq
	signal irq_mapper_receiver9_irq                                                           : std_logic;                     -- DIST2:irq -> irq_mapper:receiver9_irq
	signal irq_mapper_receiver10_irq                                                          : std_logic;                     -- DIST3:irq -> irq_mapper:receiver10_irq
	signal irq_mapper_receiver11_irq                                                          : std_logic;                     -- DIST4:irq -> irq_mapper:receiver11_irq
	signal cpu_d_irq_irq                                                                      : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:d_irq
	signal rst_controller_reset_out_reset                                                     : std_logic;                     -- rst_controller:reset_out -> [ACELEROMETRO_SPI:reset, ADC_DE0:reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                                 : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	signal rst_controller_001_reset_out_reset                                                 : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:EPCS_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal rst_controller_001_reset_out_reset_req                                             : std_logic;                     -- rst_controller_001:reset_req -> EPCS:reset_req
	signal cpu_jtag_debug_module_reset_reset                                                  : std_logic;                     -- CPU:jtag_debug_module_resetrequest -> rst_controller_001:reset_in1
	signal rst_controller_002_reset_out_reset                                                 : std_logic;                     -- rst_controller_002:reset_out -> [mm_interconnect_0:sys_pll_inclk_interface_reset_reset_bridge_in_reset_reset, sys_pll:reset]
	signal rst_controller_003_reset_out_reset                                                 : std_logic;                     -- rst_controller_003:reset_out -> [mm_interconnect_0:MOTORES_reset_reset_bridge_in_reset_reset, rst_controller_003_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                                            : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0]
	signal mm_interconnect_0_led_s1_write_ports_inv                                           : std_logic;                     -- mm_interconnect_0_led_s1_write:inv -> LED:write_n
	signal mm_interconnect_0_pwm2_s1_write_ports_inv                                          : std_logic;                     -- mm_interconnect_0_pwm2_s1_write:inv -> PWM2:write_n
	signal mm_interconnect_0_dist1_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_0_dist1_s1_write:inv -> DIST1:write_n
	signal mm_interconnect_0_dist1_s1_read_ports_inv                                          : std_logic;                     -- mm_interconnect_0_dist1_s1_read:inv -> DIST1:read_n
	signal mm_interconnect_0_gps_s1_write_ports_inv                                           : std_logic;                     -- mm_interconnect_0_gps_s1_write:inv -> GPS:write_n
	signal mm_interconnect_0_gps_s1_read_ports_inv                                            : std_logic;                     -- mm_interconnect_0_gps_s1_read:inv -> GPS:read_n
	signal mm_interconnect_0_dist3_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_0_dist3_s1_write:inv -> DIST3:write_n
	signal mm_interconnect_0_dist3_s1_read_ports_inv                                          : std_logic;                     -- mm_interconnect_0_dist3_s1_read:inv -> DIST3:read_n
	signal mm_interconnect_0_epcs_epcs_control_port_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_epcs_epcs_control_port_write:inv -> EPCS:write_n
	signal mm_interconnect_0_epcs_epcs_control_port_read_ports_inv                            : std_logic;                     -- mm_interconnect_0_epcs_epcs_control_port_read:inv -> EPCS:read_n
	signal mm_interconnect_0_xbee_s1_write_ports_inv                                          : std_logic;                     -- mm_interconnect_0_xbee_s1_write:inv -> XBEE:write_n
	signal mm_interconnect_0_xbee_s1_read_ports_inv                                           : std_logic;                     -- mm_interconnect_0_xbee_s1_read:inv -> XBEE:read_n
	signal mm_interconnect_0_sys_timer_s1_write_ports_inv                                     : std_logic;                     -- mm_interconnect_0_sys_timer_s1_write:inv -> sys_timer:write_n
	signal mm_interconnect_0_encoder_int_s1_write_ports_inv                                   : std_logic;                     -- mm_interconnect_0_encoder_int_s1_write:inv -> ENCODER_INT:write_n
	signal mm_interconnect_0_dist4_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_0_dist4_s1_write:inv -> DIST4:write_n
	signal mm_interconnect_0_dist4_s1_read_ports_inv                                          : std_logic;                     -- mm_interconnect_0_dist4_s1_read:inv -> DIST4:read_n
	signal mm_interconnect_0_data_out_i2c_s1_write_ports_inv                                  : std_logic;                     -- mm_interconnect_0_data_out_i2c_s1_write:inv -> DATA_OUT_I2C:write_n
	signal mm_interconnect_0_key_s1_write_ports_inv                                           : std_logic;                     -- mm_interconnect_0_key_s1_write:inv -> KEY:write_n
	signal mm_interconnect_0_ctrl_i2c_s1_write_ports_inv                                      : std_logic;                     -- mm_interconnect_0_ctrl_i2c_s1_write:inv -> CTRL_I2C:write_n
	signal mm_interconnect_0_motores_s1_write_ports_inv                                       : std_logic;                     -- mm_interconnect_0_motores_s1_write:inv -> MOTORES:write_n
	signal mm_interconnect_0_pwm1_s1_write_ports_inv                                          : std_logic;                     -- mm_interconnect_0_pwm1_s1_write:inv -> PWM1:write_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> SDRAM:az_wr_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                                          : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> SDRAM:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> SDRAM:az_be_n
	signal mm_interconnect_0_dist2_s1_write_ports_inv                                         : std_logic;                     -- mm_interconnect_0_dist2_s1_write:inv -> DIST2:write_n
	signal mm_interconnect_0_dist2_s1_read_ports_inv                                          : std_logic;                     -- mm_interconnect_0_dist2_s1_read:inv -> DIST2:read_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_write:inv -> JTAG:av_write_n
	signal mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv                            : std_logic;                     -- mm_interconnect_0_jtag_avalon_jtag_slave_read:inv -> JTAG:av_read_n
	signal rst_controller_reset_out_reset_ports_inv                                           : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, CTRL_I2C:reset_n, DATA_IN_I2C:reset_n, DATA_OUT_I2C:reset_n, DIST1:reset_n, DIST2:reset_n, DIST3:reset_n, DIST4:reset_n, ENCODER_INT:reset_n, ENCODER_NORMAL:reset_n, FLAG_I2C:reset_n, GPS:reset_n, JTAG:rst_n, KEY:reset_n, LED:reset_n, PWM1:reset_n, PWM2:reset_n, SDRAM:reset_n, SW:reset_n, XBEE:reset_n, sys_id:reset_n, sys_timer:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                                       : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> EPCS:reset_n
	signal rst_controller_003_reset_out_reset_ports_inv                                       : std_logic;                     -- rst_controller_003_reset_out_reset:inv -> MOTORES:reset_n

begin

	cpu : component NIOS_CPU
		port map (
			clk                                   => sys_pll_c0_clk,                                      --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,            --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                             => cpu_data_master_address,                             --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                          --                          .byteenable
			d_read                                => cpu_data_master_read,                                --                          .read
			d_readdata                            => cpu_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => cpu_data_master_write,                               --                          .write
			d_writedata                           => cpu_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                      --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                         --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                  --                          .waitrequest
			i_readdatavalid                       => cpu_instruction_master_readdatavalid,                --                          .readdatavalid
			d_irq                                 => cpu_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_cpu_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_cpu_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_cpu_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_cpu_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_cpu_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_cpu_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_cpu_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_cpu_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                 -- custom_instruction_master.readra
		);

	sys_id : component NIOS_sys_id
		port map (
			clock    => sys_pll_c0_clk,                                    --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,          --         reset.reset_n
			readdata => mm_interconnect_0_sys_id_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sys_id_control_slave_address(0)  --              .address
		);

	sdram : component NIOS_SDRAM
		port map (
			clk            => sys_pll_c0_clk,                                  --   clk.clk
			reset_n        => rst_controller_reset_out_reset_ports_inv,        -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_addr,                                      --  wire.export
			zs_ba          => sdram_ba,                                        --      .export
			zs_cas_n       => sdram_cas_n,                                     --      .export
			zs_cke         => sdram_cke,                                       --      .export
			zs_cs_n        => sdram_cs_n,                                      --      .export
			zs_dq          => sdram_dq,                                        --      .export
			zs_dqm         => sdram_dqm,                                       --      .export
			zs_ras_n       => sdram_ras_n,                                     --      .export
			zs_we_n        => sdram_we_n                                       --      .export
		);

	epcs : component NIOS_EPCS
		port map (
			clk           => sys_pll_c0_clk,                                           --               clk.clk
			reset_n       => rst_controller_001_reset_out_reset_ports_inv,             --             reset.reset_n
			reset_req     => rst_controller_001_reset_out_reset_req,                   --                  .reset_req
			address       => mm_interconnect_0_epcs_epcs_control_port_address,         -- epcs_control_port.address
			chipselect    => mm_interconnect_0_epcs_epcs_control_port_chipselect,      --                  .chipselect
			dataavailable => open,                                                     --                  .dataavailable
			endofpacket   => open,                                                     --                  .endofpacket
			read_n        => mm_interconnect_0_epcs_epcs_control_port_read_ports_inv,  --                  .read_n
			readdata      => mm_interconnect_0_epcs_epcs_control_port_readdata,        --                  .readdata
			readyfordata  => open,                                                     --                  .readyfordata
			write_n       => mm_interconnect_0_epcs_epcs_control_port_write_ports_inv, --                  .write_n
			writedata     => mm_interconnect_0_epcs_epcs_control_port_writedata,       --                  .writedata
			irq           => irq_mapper_receiver0_irq,                                 --               irq.irq
			dclk          => epcs_dclk,                                                --          external.export
			sce           => epcs_sce,                                                 --                  .export
			sdo           => epcs_sdo,                                                 --                  .export
			data0         => epcs_data0                                                --                  .export
		);

	sys_timer : component NIOS_sys_timer
		port map (
			clk        => sys_pll_c0_clk,                                 --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       -- reset.reset_n
			address    => mm_interconnect_0_sys_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_sys_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_sys_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_sys_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_sys_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                        --   irq.irq
		);

	led : component NIOS_LED
		port map (
			clk        => sys_pll_c0_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_led_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_led_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_led_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_led_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_led_s1_readdata,        --                    .readdata
			out_port   => led_export                                -- external_connection.export
		);

	sw : component NIOS_SW
		port map (
			clk      => sys_pll_c0_clk,                           --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_sw_s1_address,          --                  s1.address
			readdata => mm_interconnect_0_sw_s1_readdata,         --                    .readdata
			in_port  => sw_export                                 -- external_connection.export
		);

	key : component NIOS_KEY
		port map (
			clk        => sys_pll_c0_clk,                           --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_key_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_key_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_key_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_key_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_key_s1_readdata,        --                    .readdata
			in_port    => key_export,                               -- external_connection.export
			irq        => irq_mapper_receiver3_irq                  --                 irq.irq
		);

	jtag : component NIOS_JTAG
		port map (
			clk            => sys_pll_c0_clk,                                           --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                 --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver2_irq                                  --               irq.irq
		);

	sys_pll : component NIOS_sys_pll
		port map (
			clk       => clk_clk,                                       --       inclk_interface.clk
			reset     => rst_controller_002_reset_out_reset,            -- inclk_interface_reset.reset
			read      => mm_interconnect_0_sys_pll_pll_slave_read,      --             pll_slave.read
			write     => mm_interconnect_0_sys_pll_pll_slave_write,     --                      .write
			address   => mm_interconnect_0_sys_pll_pll_slave_address,   --                      .address
			readdata  => mm_interconnect_0_sys_pll_pll_slave_readdata,  --                      .readdata
			writedata => mm_interconnect_0_sys_pll_pll_slave_writedata, --                      .writedata
			c0        => sys_pll_c0_clk,                                --                    c0.clk
			c1        => sys_pll_c1_clk,                                --                    c1.clk
			areset    => open,                                          --        areset_conduit.export
			locked    => open,                                          --        locked_conduit.export
			phasedone => open                                           --     phasedone_conduit.export
		);

	acelerometro_spi : component NIOS_ACELEROMETRO_SPI
		port map (
			clk           => sys_pll_c0_clk,                                                                       --                         clock_reset.clk
			reset         => rst_controller_reset_out_reset,                                                       --                   clock_reset_reset.reset
			address       => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_address(0),    -- avalon_accelerometer_spi_mode_slave.address
			byteenable    => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_byteenable(0), --                                    .byteenable
			read          => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_read,          --                                    .read
			write         => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_write,         --                                    .write
			writedata     => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_writedata,     --                                    .writedata
			readdata      => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_readdata,      --                                    .readdata
			waitrequest   => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_waitrequest,   --                                    .waitrequest
			irq           => irq_mapper_receiver5_irq,                                                             --                           interrupt.irq
			I2C_SDAT      => acelerometro_spi_I2C_SDAT,                                                            --                  external_interface.export
			I2C_SCLK      => acelerometro_spi_I2C_SCLK,                                                            --                                    .export
			G_SENSOR_CS_N => acelerometro_spi_G_SENSOR_CS_N,                                                       --                                    .export
			G_SENSOR_INT  => acelerometro_spi_G_SENSOR_INT                                                         --                                    .export
		);

	adc_de0 : component NIOS_ADC_DE0
		port map (
			clock       => sys_pll_c0_clk,                                  --                clk.clk
			reset       => rst_controller_reset_out_reset,                  --              reset.reset
			write       => mm_interconnect_0_adc_de0_adc_slave_write,       --          adc_slave.write
			readdata    => mm_interconnect_0_adc_de0_adc_slave_readdata,    --                   .readdata
			writedata   => mm_interconnect_0_adc_de0_adc_slave_writedata,   --                   .writedata
			address     => mm_interconnect_0_adc_de0_adc_slave_address,     --                   .address
			waitrequest => mm_interconnect_0_adc_de0_adc_slave_waitrequest, --                   .waitrequest
			read        => mm_interconnect_0_adc_de0_adc_slave_read,        --                   .read
			adc_sclk    => adc_sclk,                                        -- external_interface.export
			adc_cs_n    => adc_cs_n,                                        --                   .export
			adc_dout    => adc_dout,                                        --                   .export
			adc_din     => adc_din                                          --                   .export
		);

	encoder_int : component NIOS_ENCODER_INT
		port map (
			clk        => sys_pll_c0_clk,                                   --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,         --               reset.reset_n
			address    => mm_interconnect_0_encoder_int_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_encoder_int_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_encoder_int_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_encoder_int_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_encoder_int_s1_readdata,        --                    .readdata
			in_port    => encoder_int_export,                               -- external_connection.export
			irq        => irq_mapper_receiver4_irq                          --                 irq.irq
		);

	encoder_normal : component NIOS_SW
		port map (
			clk      => sys_pll_c0_clk,                               --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address  => mm_interconnect_0_encoder_normal_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_encoder_normal_s1_readdata, --                    .readdata
			in_port  => encoder_normal_export                         -- external_connection.export
		);

	motores : component NIOS_MOTORES
		port map (
			clk        => sys_pll_c1_clk,                               --                 clk.clk
			reset_n    => rst_controller_003_reset_out_reset_ports_inv, --               reset.reset_n
			address    => mm_interconnect_0_motores_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_motores_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_motores_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_motores_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_motores_s1_readdata,        --                    .readdata
			out_port   => motores_export                                -- external_connection.export
		);

	pwm1 : component NIOS_LED
		port map (
			clk        => sys_pll_c0_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_pwm1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm1_s1_readdata,        --                    .readdata
			out_port   => pwm1_export                                -- external_connection.export
		);

	pwm2 : component NIOS_LED
		port map (
			clk        => sys_pll_c0_clk,                            --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address    => mm_interconnect_0_pwm2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pwm2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pwm2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pwm2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pwm2_s1_readdata,        --                    .readdata
			out_port   => pwm2_export                                -- external_connection.export
		);

	ctrl_i2c : component NIOS_CTRL_I2C
		port map (
			clk        => sys_pll_c0_clk,                                --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_ctrl_i2c_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_ctrl_i2c_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_ctrl_i2c_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_ctrl_i2c_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_ctrl_i2c_s1_readdata,        --                    .readdata
			out_port   => ctrl_i2c_export                                -- external_connection.export
		);

	data_out_i2c : component NIOS_LED
		port map (
			clk        => sys_pll_c0_clk,                                    --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,          --               reset.reset_n
			address    => mm_interconnect_0_data_out_i2c_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_data_out_i2c_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_data_out_i2c_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_data_out_i2c_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_data_out_i2c_s1_readdata,        --                    .readdata
			out_port   => data_out_i2c_export                                -- external_connection.export
		);

	data_in_i2c : component NIOS_DATA_IN_I2C
		port map (
			clk      => sys_pll_c0_clk,                            --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => mm_interconnect_0_data_in_i2c_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_data_in_i2c_s1_readdata, --                    .readdata
			in_port  => data_in_i2c_export                         -- external_connection.export
		);

	flag_i2c : component NIOS_FLAG_I2C
		port map (
			clk      => sys_pll_c0_clk,                           --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_flag_i2c_s1_address,    --                  s1.address
			readdata => mm_interconnect_0_flag_i2c_s1_readdata,   --                    .readdata
			in_port  => flag_i2c_export                           -- external_connection.export
		);

	gps : component NIOS_GPS
		port map (
			clk           => sys_pll_c0_clk,                           --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address       => mm_interconnect_0_gps_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_gps_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_gps_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_gps_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_gps_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_gps_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_gps_s1_readdata,        --                    .readdata
			dataavailable => open,                                     --                    .dataavailable
			readyfordata  => open,                                     --                    .readyfordata
			rxd           => gps_rxd,                                  -- external_connection.export
			txd           => gps_txd,                                  --                    .export
			irq           => irq_mapper_receiver6_irq                  --                 irq.irq
		);

	xbee : component NIOS_GPS
		port map (
			clk           => sys_pll_c0_clk,                            --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address       => mm_interconnect_0_xbee_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_xbee_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_xbee_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_xbee_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_xbee_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_xbee_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_xbee_s1_readdata,        --                    .readdata
			dataavailable => open,                                      --                    .dataavailable
			readyfordata  => open,                                      --                    .readyfordata
			rxd           => xbee_rxd,                                  -- external_connection.export
			txd           => xbee_txd,                                  --                    .export
			irq           => irq_mapper_receiver7_irq                   --                 irq.irq
		);

	dist1 : component NIOS_GPS
		port map (
			clk           => sys_pll_c0_clk,                             --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address       => mm_interconnect_0_dist1_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_dist1_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_dist1_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_dist1_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_dist1_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_dist1_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_dist1_s1_readdata,        --                    .readdata
			dataavailable => open,                                       --                    .dataavailable
			readyfordata  => open,                                       --                    .readyfordata
			rxd           => dist1_rxd,                                  -- external_connection.export
			txd           => dist1_txd,                                  --                    .export
			irq           => irq_mapper_receiver8_irq                    --                 irq.irq
		);

	dist2 : component NIOS_GPS
		port map (
			clk           => sys_pll_c0_clk,                             --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address       => mm_interconnect_0_dist2_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_dist2_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_dist2_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_dist2_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_dist2_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_dist2_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_dist2_s1_readdata,        --                    .readdata
			dataavailable => open,                                       --                    .dataavailable
			readyfordata  => open,                                       --                    .readyfordata
			rxd           => dist2_rxd,                                  -- external_connection.export
			txd           => dist2_txd,                                  --                    .export
			irq           => irq_mapper_receiver9_irq                    --                 irq.irq
		);

	dist3 : component NIOS_GPS
		port map (
			clk           => sys_pll_c0_clk,                             --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address       => mm_interconnect_0_dist3_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_dist3_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_dist3_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_dist3_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_dist3_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_dist3_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_dist3_s1_readdata,        --                    .readdata
			dataavailable => open,                                       --                    .dataavailable
			readyfordata  => open,                                       --                    .readyfordata
			rxd           => dist3_rxd,                                  -- external_connection.export
			txd           => dist3_txd,                                  --                    .export
			irq           => irq_mapper_receiver10_irq                   --                 irq.irq
		);

	dist4 : component NIOS_GPS
		port map (
			clk           => sys_pll_c0_clk,                             --                 clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,   --               reset.reset_n
			address       => mm_interconnect_0_dist4_s1_address,         --                  s1.address
			begintransfer => mm_interconnect_0_dist4_s1_begintransfer,   --                    .begintransfer
			chipselect    => mm_interconnect_0_dist4_s1_chipselect,      --                    .chipselect
			read_n        => mm_interconnect_0_dist4_s1_read_ports_inv,  --                    .read_n
			write_n       => mm_interconnect_0_dist4_s1_write_ports_inv, --                    .write_n
			writedata     => mm_interconnect_0_dist4_s1_writedata,       --                    .writedata
			readdata      => mm_interconnect_0_dist4_s1_readdata,        --                    .readdata
			dataavailable => open,                                       --                    .dataavailable
			readyfordata  => open,                                       --                    .readyfordata
			rxd           => dist4_rxd,                                  -- external_connection.export
			txd           => dist4_txd,                                  --                    .export
			irq           => irq_mapper_receiver11_irq                   --                 irq.irq
		);

	mm_interconnect_0 : component NIOS_mm_interconnect_0
		port map (
			clk_50_clk_clk                                                   => clk_clk,                                                                            --                                           clk_50_clk.clk
			ram_clk_clk_clk                                                  => sys_pll_c1_clk,                                                                     --                                          ram_clk_clk.clk
			sys_clk_clk_clk                                                  => sys_pll_c0_clk,                                                                     --                                          sys_clk_clk.clk
			CPU_reset_n_reset_bridge_in_reset_reset                          => rst_controller_reset_out_reset,                                                     --                    CPU_reset_n_reset_bridge_in_reset.reset
			EPCS_reset_reset_bridge_in_reset_reset                           => rst_controller_001_reset_out_reset,                                                 --                     EPCS_reset_reset_bridge_in_reset.reset
			MOTORES_reset_reset_bridge_in_reset_reset                        => rst_controller_003_reset_out_reset,                                                 --                  MOTORES_reset_reset_bridge_in_reset.reset
			sys_pll_inclk_interface_reset_reset_bridge_in_reset_reset        => rst_controller_002_reset_out_reset,                                                 --  sys_pll_inclk_interface_reset_reset_bridge_in_reset.reset
			CPU_data_master_address                                          => cpu_data_master_address,                                                            --                                      CPU_data_master.address
			CPU_data_master_waitrequest                                      => cpu_data_master_waitrequest,                                                        --                                                     .waitrequest
			CPU_data_master_byteenable                                       => cpu_data_master_byteenable,                                                         --                                                     .byteenable
			CPU_data_master_read                                             => cpu_data_master_read,                                                               --                                                     .read
			CPU_data_master_readdata                                         => cpu_data_master_readdata,                                                           --                                                     .readdata
			CPU_data_master_write                                            => cpu_data_master_write,                                                              --                                                     .write
			CPU_data_master_writedata                                        => cpu_data_master_writedata,                                                          --                                                     .writedata
			CPU_data_master_debugaccess                                      => cpu_data_master_debugaccess,                                                        --                                                     .debugaccess
			CPU_instruction_master_address                                   => cpu_instruction_master_address,                                                     --                               CPU_instruction_master.address
			CPU_instruction_master_waitrequest                               => cpu_instruction_master_waitrequest,                                                 --                                                     .waitrequest
			CPU_instruction_master_read                                      => cpu_instruction_master_read,                                                        --                                                     .read
			CPU_instruction_master_readdata                                  => cpu_instruction_master_readdata,                                                    --                                                     .readdata
			CPU_instruction_master_readdatavalid                             => cpu_instruction_master_readdatavalid,                                               --                                                     .readdatavalid
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_address     => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_address,     -- ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave.address
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_write       => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_write,       --                                                     .write
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_read        => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_read,        --                                                     .read
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_readdata    => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_readdata,    --                                                     .readdata
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_writedata   => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_writedata,   --                                                     .writedata
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_byteenable  => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_byteenable,  --                                                     .byteenable
			ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_waitrequest => mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_waitrequest, --                                                     .waitrequest
			ADC_DE0_adc_slave_address                                        => mm_interconnect_0_adc_de0_adc_slave_address,                                        --                                    ADC_DE0_adc_slave.address
			ADC_DE0_adc_slave_write                                          => mm_interconnect_0_adc_de0_adc_slave_write,                                          --                                                     .write
			ADC_DE0_adc_slave_read                                           => mm_interconnect_0_adc_de0_adc_slave_read,                                           --                                                     .read
			ADC_DE0_adc_slave_readdata                                       => mm_interconnect_0_adc_de0_adc_slave_readdata,                                       --                                                     .readdata
			ADC_DE0_adc_slave_writedata                                      => mm_interconnect_0_adc_de0_adc_slave_writedata,                                      --                                                     .writedata
			ADC_DE0_adc_slave_waitrequest                                    => mm_interconnect_0_adc_de0_adc_slave_waitrequest,                                    --                                                     .waitrequest
			CPU_jtag_debug_module_address                                    => mm_interconnect_0_cpu_jtag_debug_module_address,                                    --                                CPU_jtag_debug_module.address
			CPU_jtag_debug_module_write                                      => mm_interconnect_0_cpu_jtag_debug_module_write,                                      --                                                     .write
			CPU_jtag_debug_module_read                                       => mm_interconnect_0_cpu_jtag_debug_module_read,                                       --                                                     .read
			CPU_jtag_debug_module_readdata                                   => mm_interconnect_0_cpu_jtag_debug_module_readdata,                                   --                                                     .readdata
			CPU_jtag_debug_module_writedata                                  => mm_interconnect_0_cpu_jtag_debug_module_writedata,                                  --                                                     .writedata
			CPU_jtag_debug_module_byteenable                                 => mm_interconnect_0_cpu_jtag_debug_module_byteenable,                                 --                                                     .byteenable
			CPU_jtag_debug_module_waitrequest                                => mm_interconnect_0_cpu_jtag_debug_module_waitrequest,                                --                                                     .waitrequest
			CPU_jtag_debug_module_debugaccess                                => mm_interconnect_0_cpu_jtag_debug_module_debugaccess,                                --                                                     .debugaccess
			CTRL_I2C_s1_address                                              => mm_interconnect_0_ctrl_i2c_s1_address,                                              --                                          CTRL_I2C_s1.address
			CTRL_I2C_s1_write                                                => mm_interconnect_0_ctrl_i2c_s1_write,                                                --                                                     .write
			CTRL_I2C_s1_readdata                                             => mm_interconnect_0_ctrl_i2c_s1_readdata,                                             --                                                     .readdata
			CTRL_I2C_s1_writedata                                            => mm_interconnect_0_ctrl_i2c_s1_writedata,                                            --                                                     .writedata
			CTRL_I2C_s1_chipselect                                           => mm_interconnect_0_ctrl_i2c_s1_chipselect,                                           --                                                     .chipselect
			DATA_IN_I2C_s1_address                                           => mm_interconnect_0_data_in_i2c_s1_address,                                           --                                       DATA_IN_I2C_s1.address
			DATA_IN_I2C_s1_readdata                                          => mm_interconnect_0_data_in_i2c_s1_readdata,                                          --                                                     .readdata
			DATA_OUT_I2C_s1_address                                          => mm_interconnect_0_data_out_i2c_s1_address,                                          --                                      DATA_OUT_I2C_s1.address
			DATA_OUT_I2C_s1_write                                            => mm_interconnect_0_data_out_i2c_s1_write,                                            --                                                     .write
			DATA_OUT_I2C_s1_readdata                                         => mm_interconnect_0_data_out_i2c_s1_readdata,                                         --                                                     .readdata
			DATA_OUT_I2C_s1_writedata                                        => mm_interconnect_0_data_out_i2c_s1_writedata,                                        --                                                     .writedata
			DATA_OUT_I2C_s1_chipselect                                       => mm_interconnect_0_data_out_i2c_s1_chipselect,                                       --                                                     .chipselect
			DIST1_s1_address                                                 => mm_interconnect_0_dist1_s1_address,                                                 --                                             DIST1_s1.address
			DIST1_s1_write                                                   => mm_interconnect_0_dist1_s1_write,                                                   --                                                     .write
			DIST1_s1_read                                                    => mm_interconnect_0_dist1_s1_read,                                                    --                                                     .read
			DIST1_s1_readdata                                                => mm_interconnect_0_dist1_s1_readdata,                                                --                                                     .readdata
			DIST1_s1_writedata                                               => mm_interconnect_0_dist1_s1_writedata,                                               --                                                     .writedata
			DIST1_s1_begintransfer                                           => mm_interconnect_0_dist1_s1_begintransfer,                                           --                                                     .begintransfer
			DIST1_s1_chipselect                                              => mm_interconnect_0_dist1_s1_chipselect,                                              --                                                     .chipselect
			DIST2_s1_address                                                 => mm_interconnect_0_dist2_s1_address,                                                 --                                             DIST2_s1.address
			DIST2_s1_write                                                   => mm_interconnect_0_dist2_s1_write,                                                   --                                                     .write
			DIST2_s1_read                                                    => mm_interconnect_0_dist2_s1_read,                                                    --                                                     .read
			DIST2_s1_readdata                                                => mm_interconnect_0_dist2_s1_readdata,                                                --                                                     .readdata
			DIST2_s1_writedata                                               => mm_interconnect_0_dist2_s1_writedata,                                               --                                                     .writedata
			DIST2_s1_begintransfer                                           => mm_interconnect_0_dist2_s1_begintransfer,                                           --                                                     .begintransfer
			DIST2_s1_chipselect                                              => mm_interconnect_0_dist2_s1_chipselect,                                              --                                                     .chipselect
			DIST3_s1_address                                                 => mm_interconnect_0_dist3_s1_address,                                                 --                                             DIST3_s1.address
			DIST3_s1_write                                                   => mm_interconnect_0_dist3_s1_write,                                                   --                                                     .write
			DIST3_s1_read                                                    => mm_interconnect_0_dist3_s1_read,                                                    --                                                     .read
			DIST3_s1_readdata                                                => mm_interconnect_0_dist3_s1_readdata,                                                --                                                     .readdata
			DIST3_s1_writedata                                               => mm_interconnect_0_dist3_s1_writedata,                                               --                                                     .writedata
			DIST3_s1_begintransfer                                           => mm_interconnect_0_dist3_s1_begintransfer,                                           --                                                     .begintransfer
			DIST3_s1_chipselect                                              => mm_interconnect_0_dist3_s1_chipselect,                                              --                                                     .chipselect
			DIST4_s1_address                                                 => mm_interconnect_0_dist4_s1_address,                                                 --                                             DIST4_s1.address
			DIST4_s1_write                                                   => mm_interconnect_0_dist4_s1_write,                                                   --                                                     .write
			DIST4_s1_read                                                    => mm_interconnect_0_dist4_s1_read,                                                    --                                                     .read
			DIST4_s1_readdata                                                => mm_interconnect_0_dist4_s1_readdata,                                                --                                                     .readdata
			DIST4_s1_writedata                                               => mm_interconnect_0_dist4_s1_writedata,                                               --                                                     .writedata
			DIST4_s1_begintransfer                                           => mm_interconnect_0_dist4_s1_begintransfer,                                           --                                                     .begintransfer
			DIST4_s1_chipselect                                              => mm_interconnect_0_dist4_s1_chipselect,                                              --                                                     .chipselect
			ENCODER_INT_s1_address                                           => mm_interconnect_0_encoder_int_s1_address,                                           --                                       ENCODER_INT_s1.address
			ENCODER_INT_s1_write                                             => mm_interconnect_0_encoder_int_s1_write,                                             --                                                     .write
			ENCODER_INT_s1_readdata                                          => mm_interconnect_0_encoder_int_s1_readdata,                                          --                                                     .readdata
			ENCODER_INT_s1_writedata                                         => mm_interconnect_0_encoder_int_s1_writedata,                                         --                                                     .writedata
			ENCODER_INT_s1_chipselect                                        => mm_interconnect_0_encoder_int_s1_chipselect,                                        --                                                     .chipselect
			ENCODER_NORMAL_s1_address                                        => mm_interconnect_0_encoder_normal_s1_address,                                        --                                    ENCODER_NORMAL_s1.address
			ENCODER_NORMAL_s1_readdata                                       => mm_interconnect_0_encoder_normal_s1_readdata,                                       --                                                     .readdata
			EPCS_epcs_control_port_address                                   => mm_interconnect_0_epcs_epcs_control_port_address,                                   --                               EPCS_epcs_control_port.address
			EPCS_epcs_control_port_write                                     => mm_interconnect_0_epcs_epcs_control_port_write,                                     --                                                     .write
			EPCS_epcs_control_port_read                                      => mm_interconnect_0_epcs_epcs_control_port_read,                                      --                                                     .read
			EPCS_epcs_control_port_readdata                                  => mm_interconnect_0_epcs_epcs_control_port_readdata,                                  --                                                     .readdata
			EPCS_epcs_control_port_writedata                                 => mm_interconnect_0_epcs_epcs_control_port_writedata,                                 --                                                     .writedata
			EPCS_epcs_control_port_chipselect                                => mm_interconnect_0_epcs_epcs_control_port_chipselect,                                --                                                     .chipselect
			FLAG_I2C_s1_address                                              => mm_interconnect_0_flag_i2c_s1_address,                                              --                                          FLAG_I2C_s1.address
			FLAG_I2C_s1_readdata                                             => mm_interconnect_0_flag_i2c_s1_readdata,                                             --                                                     .readdata
			GPS_s1_address                                                   => mm_interconnect_0_gps_s1_address,                                                   --                                               GPS_s1.address
			GPS_s1_write                                                     => mm_interconnect_0_gps_s1_write,                                                     --                                                     .write
			GPS_s1_read                                                      => mm_interconnect_0_gps_s1_read,                                                      --                                                     .read
			GPS_s1_readdata                                                  => mm_interconnect_0_gps_s1_readdata,                                                  --                                                     .readdata
			GPS_s1_writedata                                                 => mm_interconnect_0_gps_s1_writedata,                                                 --                                                     .writedata
			GPS_s1_begintransfer                                             => mm_interconnect_0_gps_s1_begintransfer,                                             --                                                     .begintransfer
			GPS_s1_chipselect                                                => mm_interconnect_0_gps_s1_chipselect,                                                --                                                     .chipselect
			JTAG_avalon_jtag_slave_address                                   => mm_interconnect_0_jtag_avalon_jtag_slave_address,                                   --                               JTAG_avalon_jtag_slave.address
			JTAG_avalon_jtag_slave_write                                     => mm_interconnect_0_jtag_avalon_jtag_slave_write,                                     --                                                     .write
			JTAG_avalon_jtag_slave_read                                      => mm_interconnect_0_jtag_avalon_jtag_slave_read,                                      --                                                     .read
			JTAG_avalon_jtag_slave_readdata                                  => mm_interconnect_0_jtag_avalon_jtag_slave_readdata,                                  --                                                     .readdata
			JTAG_avalon_jtag_slave_writedata                                 => mm_interconnect_0_jtag_avalon_jtag_slave_writedata,                                 --                                                     .writedata
			JTAG_avalon_jtag_slave_waitrequest                               => mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest,                               --                                                     .waitrequest
			JTAG_avalon_jtag_slave_chipselect                                => mm_interconnect_0_jtag_avalon_jtag_slave_chipselect,                                --                                                     .chipselect
			KEY_s1_address                                                   => mm_interconnect_0_key_s1_address,                                                   --                                               KEY_s1.address
			KEY_s1_write                                                     => mm_interconnect_0_key_s1_write,                                                     --                                                     .write
			KEY_s1_readdata                                                  => mm_interconnect_0_key_s1_readdata,                                                  --                                                     .readdata
			KEY_s1_writedata                                                 => mm_interconnect_0_key_s1_writedata,                                                 --                                                     .writedata
			KEY_s1_chipselect                                                => mm_interconnect_0_key_s1_chipselect,                                                --                                                     .chipselect
			LED_s1_address                                                   => mm_interconnect_0_led_s1_address,                                                   --                                               LED_s1.address
			LED_s1_write                                                     => mm_interconnect_0_led_s1_write,                                                     --                                                     .write
			LED_s1_readdata                                                  => mm_interconnect_0_led_s1_readdata,                                                  --                                                     .readdata
			LED_s1_writedata                                                 => mm_interconnect_0_led_s1_writedata,                                                 --                                                     .writedata
			LED_s1_chipselect                                                => mm_interconnect_0_led_s1_chipselect,                                                --                                                     .chipselect
			MOTORES_s1_address                                               => mm_interconnect_0_motores_s1_address,                                               --                                           MOTORES_s1.address
			MOTORES_s1_write                                                 => mm_interconnect_0_motores_s1_write,                                                 --                                                     .write
			MOTORES_s1_readdata                                              => mm_interconnect_0_motores_s1_readdata,                                              --                                                     .readdata
			MOTORES_s1_writedata                                             => mm_interconnect_0_motores_s1_writedata,                                             --                                                     .writedata
			MOTORES_s1_chipselect                                            => mm_interconnect_0_motores_s1_chipselect,                                            --                                                     .chipselect
			PWM1_s1_address                                                  => mm_interconnect_0_pwm1_s1_address,                                                  --                                              PWM1_s1.address
			PWM1_s1_write                                                    => mm_interconnect_0_pwm1_s1_write,                                                    --                                                     .write
			PWM1_s1_readdata                                                 => mm_interconnect_0_pwm1_s1_readdata,                                                 --                                                     .readdata
			PWM1_s1_writedata                                                => mm_interconnect_0_pwm1_s1_writedata,                                                --                                                     .writedata
			PWM1_s1_chipselect                                               => mm_interconnect_0_pwm1_s1_chipselect,                                               --                                                     .chipselect
			PWM2_s1_address                                                  => mm_interconnect_0_pwm2_s1_address,                                                  --                                              PWM2_s1.address
			PWM2_s1_write                                                    => mm_interconnect_0_pwm2_s1_write,                                                    --                                                     .write
			PWM2_s1_readdata                                                 => mm_interconnect_0_pwm2_s1_readdata,                                                 --                                                     .readdata
			PWM2_s1_writedata                                                => mm_interconnect_0_pwm2_s1_writedata,                                                --                                                     .writedata
			PWM2_s1_chipselect                                               => mm_interconnect_0_pwm2_s1_chipselect,                                               --                                                     .chipselect
			SDRAM_s1_address                                                 => mm_interconnect_0_sdram_s1_address,                                                 --                                             SDRAM_s1.address
			SDRAM_s1_write                                                   => mm_interconnect_0_sdram_s1_write,                                                   --                                                     .write
			SDRAM_s1_read                                                    => mm_interconnect_0_sdram_s1_read,                                                    --                                                     .read
			SDRAM_s1_readdata                                                => mm_interconnect_0_sdram_s1_readdata,                                                --                                                     .readdata
			SDRAM_s1_writedata                                               => mm_interconnect_0_sdram_s1_writedata,                                               --                                                     .writedata
			SDRAM_s1_byteenable                                              => mm_interconnect_0_sdram_s1_byteenable,                                              --                                                     .byteenable
			SDRAM_s1_readdatavalid                                           => mm_interconnect_0_sdram_s1_readdatavalid,                                           --                                                     .readdatavalid
			SDRAM_s1_waitrequest                                             => mm_interconnect_0_sdram_s1_waitrequest,                                             --                                                     .waitrequest
			SDRAM_s1_chipselect                                              => mm_interconnect_0_sdram_s1_chipselect,                                              --                                                     .chipselect
			SW_s1_address                                                    => mm_interconnect_0_sw_s1_address,                                                    --                                                SW_s1.address
			SW_s1_readdata                                                   => mm_interconnect_0_sw_s1_readdata,                                                   --                                                     .readdata
			sys_id_control_slave_address                                     => mm_interconnect_0_sys_id_control_slave_address,                                     --                                 sys_id_control_slave.address
			sys_id_control_slave_readdata                                    => mm_interconnect_0_sys_id_control_slave_readdata,                                    --                                                     .readdata
			sys_pll_pll_slave_address                                        => mm_interconnect_0_sys_pll_pll_slave_address,                                        --                                    sys_pll_pll_slave.address
			sys_pll_pll_slave_write                                          => mm_interconnect_0_sys_pll_pll_slave_write,                                          --                                                     .write
			sys_pll_pll_slave_read                                           => mm_interconnect_0_sys_pll_pll_slave_read,                                           --                                                     .read
			sys_pll_pll_slave_readdata                                       => mm_interconnect_0_sys_pll_pll_slave_readdata,                                       --                                                     .readdata
			sys_pll_pll_slave_writedata                                      => mm_interconnect_0_sys_pll_pll_slave_writedata,                                      --                                                     .writedata
			sys_timer_s1_address                                             => mm_interconnect_0_sys_timer_s1_address,                                             --                                         sys_timer_s1.address
			sys_timer_s1_write                                               => mm_interconnect_0_sys_timer_s1_write,                                               --                                                     .write
			sys_timer_s1_readdata                                            => mm_interconnect_0_sys_timer_s1_readdata,                                            --                                                     .readdata
			sys_timer_s1_writedata                                           => mm_interconnect_0_sys_timer_s1_writedata,                                           --                                                     .writedata
			sys_timer_s1_chipselect                                          => mm_interconnect_0_sys_timer_s1_chipselect,                                          --                                                     .chipselect
			XBEE_s1_address                                                  => mm_interconnect_0_xbee_s1_address,                                                  --                                              XBEE_s1.address
			XBEE_s1_write                                                    => mm_interconnect_0_xbee_s1_write,                                                    --                                                     .write
			XBEE_s1_read                                                     => mm_interconnect_0_xbee_s1_read,                                                     --                                                     .read
			XBEE_s1_readdata                                                 => mm_interconnect_0_xbee_s1_readdata,                                                 --                                                     .readdata
			XBEE_s1_writedata                                                => mm_interconnect_0_xbee_s1_writedata,                                                --                                                     .writedata
			XBEE_s1_begintransfer                                            => mm_interconnect_0_xbee_s1_begintransfer,                                            --                                                     .begintransfer
			XBEE_s1_chipselect                                               => mm_interconnect_0_xbee_s1_chipselect                                                --                                                     .chipselect
		);

	irq_mapper : component NIOS_irq_mapper
		port map (
			clk            => sys_pll_c0_clk,                 --        clk.clk
			reset          => rst_controller_reset_out_reset, --  clk_reset.reset
			receiver0_irq  => irq_mapper_receiver0_irq,       --  receiver0.irq
			receiver1_irq  => irq_mapper_receiver1_irq,       --  receiver1.irq
			receiver2_irq  => irq_mapper_receiver2_irq,       --  receiver2.irq
			receiver3_irq  => irq_mapper_receiver3_irq,       --  receiver3.irq
			receiver4_irq  => irq_mapper_receiver4_irq,       --  receiver4.irq
			receiver5_irq  => irq_mapper_receiver5_irq,       --  receiver5.irq
			receiver6_irq  => irq_mapper_receiver6_irq,       --  receiver6.irq
			receiver7_irq  => irq_mapper_receiver7_irq,       --  receiver7.irq
			receiver8_irq  => irq_mapper_receiver8_irq,       --  receiver8.irq
			receiver9_irq  => irq_mapper_receiver9_irq,       --  receiver9.irq
			receiver10_irq => irq_mapper_receiver10_irq,      -- receiver10.irq
			receiver11_irq => irq_mapper_receiver11_irq,      -- receiver11.irq
			sender_irq     => cpu_d_irq_irq                   --     sender.irq
		);

	rst_controller : component nios_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => sys_pll_c0_clk,                     --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component nios_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => cpu_jtag_debug_module_reset_reset,      -- reset_in1.reset
			clk            => sys_pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_001_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_002 : component nios_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_002_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_003 : component nios_rst_controller_002
		generic map (
			NUM_RESET_INPUTS          => 1,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			clk            => sys_pll_c1_clk,                     --       clk.clk
			reset_out      => rst_controller_003_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_in1      => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_led_s1_write_ports_inv <= not mm_interconnect_0_led_s1_write;

	mm_interconnect_0_pwm2_s1_write_ports_inv <= not mm_interconnect_0_pwm2_s1_write;

	mm_interconnect_0_dist1_s1_write_ports_inv <= not mm_interconnect_0_dist1_s1_write;

	mm_interconnect_0_dist1_s1_read_ports_inv <= not mm_interconnect_0_dist1_s1_read;

	mm_interconnect_0_gps_s1_write_ports_inv <= not mm_interconnect_0_gps_s1_write;

	mm_interconnect_0_gps_s1_read_ports_inv <= not mm_interconnect_0_gps_s1_read;

	mm_interconnect_0_dist3_s1_write_ports_inv <= not mm_interconnect_0_dist3_s1_write;

	mm_interconnect_0_dist3_s1_read_ports_inv <= not mm_interconnect_0_dist3_s1_read;

	mm_interconnect_0_epcs_epcs_control_port_write_ports_inv <= not mm_interconnect_0_epcs_epcs_control_port_write;

	mm_interconnect_0_epcs_epcs_control_port_read_ports_inv <= not mm_interconnect_0_epcs_epcs_control_port_read;

	mm_interconnect_0_xbee_s1_write_ports_inv <= not mm_interconnect_0_xbee_s1_write;

	mm_interconnect_0_xbee_s1_read_ports_inv <= not mm_interconnect_0_xbee_s1_read;

	mm_interconnect_0_sys_timer_s1_write_ports_inv <= not mm_interconnect_0_sys_timer_s1_write;

	mm_interconnect_0_encoder_int_s1_write_ports_inv <= not mm_interconnect_0_encoder_int_s1_write;

	mm_interconnect_0_dist4_s1_write_ports_inv <= not mm_interconnect_0_dist4_s1_write;

	mm_interconnect_0_dist4_s1_read_ports_inv <= not mm_interconnect_0_dist4_s1_read;

	mm_interconnect_0_data_out_i2c_s1_write_ports_inv <= not mm_interconnect_0_data_out_i2c_s1_write;

	mm_interconnect_0_key_s1_write_ports_inv <= not mm_interconnect_0_key_s1_write;

	mm_interconnect_0_ctrl_i2c_s1_write_ports_inv <= not mm_interconnect_0_ctrl_i2c_s1_write;

	mm_interconnect_0_motores_s1_write_ports_inv <= not mm_interconnect_0_motores_s1_write;

	mm_interconnect_0_pwm1_s1_write_ports_inv <= not mm_interconnect_0_pwm1_s1_write;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_dist2_s1_write_ports_inv <= not mm_interconnect_0_dist2_s1_write;

	mm_interconnect_0_dist2_s1_read_ports_inv <= not mm_interconnect_0_dist2_s1_read;

	mm_interconnect_0_jtag_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_avalon_jtag_slave_read;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

	rst_controller_003_reset_out_reset_ports_inv <= not rst_controller_003_reset_out_reset;

end architecture rtl; -- of NIOS
