// NIOS.v

// Generated using ACDS version 13.1 182 at 2019.09.20.11:23:32

`timescale 1 ps / 1 ps
module NIOS (
		input  wire        clk_clk,                        //              clk.clk
		input  wire        reset_reset_n,                  //            reset.reset_n
		output wire [12:0] sdram_addr,                     //            sdram.addr
		output wire [1:0]  sdram_ba,                       //                 .ba
		output wire        sdram_cas_n,                    //                 .cas_n
		output wire        sdram_cke,                      //                 .cke
		output wire        sdram_cs_n,                     //                 .cs_n
		inout  wire [15:0] sdram_dq,                       //                 .dq
		output wire [1:0]  sdram_dqm,                      //                 .dqm
		output wire        sdram_ras_n,                    //                 .ras_n
		output wire        sdram_we_n,                     //                 .we_n
		output wire        epcs_dclk,                      //             epcs.dclk
		output wire        epcs_sce,                       //                 .sce
		output wire        epcs_sdo,                       //                 .sdo
		input  wire        epcs_data0,                     //                 .data0
		output wire [7:0]  led_export,                     //              led.export
		input  wire [3:0]  sw_export,                      //               sw.export
		input  wire [1:0]  key_export,                     //              key.export
		output wire        ram_clk_clk,                    //          ram_clk.clk
		inout  wire        acelerometro_spi_I2C_SDAT,      // acelerometro_spi.I2C_SDAT
		output wire        acelerometro_spi_I2C_SCLK,      //                 .I2C_SCLK
		output wire        acelerometro_spi_G_SENSOR_CS_N, //                 .G_SENSOR_CS_N
		input  wire        acelerometro_spi_G_SENSOR_INT,  //                 .G_SENSOR_INT
		output wire        adc_sclk,                       //              adc.sclk
		output wire        adc_cs_n,                       //                 .cs_n
		input  wire        adc_dout,                       //                 .dout
		output wire        adc_din,                        //                 .din
		input  wire [3:0]  encoder_int_export,             //      encoder_int.export
		input  wire [3:0]  encoder_normal_export,          //   encoder_normal.export
		output wire [5:0]  motores_export,                 //          motores.export
		output wire [7:0]  pwm1_export,                    //             pwm1.export
		output wire [7:0]  pwm2_export,                    //             pwm2.export
		output wire [6:0]  ctrl_i2c_export,                //         ctrl_i2c.export
		output wire [7:0]  data_out_i2c_export,            //     data_out_i2c.export
		input  wire [7:0]  data_in_i2c_export,             //      data_in_i2c.export
		input  wire [1:0]  flag_i2c_export,                //         flag_i2c.export
		input  wire        gps_rxd,                        //              gps.rxd
		output wire        gps_txd,                        //                 .txd
		input  wire        xbee_rxd,                       //             xbee.rxd
		output wire        xbee_txd,                       //                 .txd
		input  wire        dist1_rxd,                      //            dist1.rxd
		output wire        dist1_txd,                      //                 .txd
		input  wire        dist2_rxd,                      //            dist2.rxd
		output wire        dist2_txd,                      //                 .txd
		input  wire        dist3_rxd,                      //            dist3.rxd
		output wire        dist3_txd,                      //                 .txd
		input  wire        dist4_rxd,                      //            dist4.rxd
		output wire        dist4_txd,                      //                 .txd
		input  wire        dist5_rxd,                      //            dist5.rxd
		output wire        dist5_txd,                      //                 .txd
		input  wire        dist6_rxd,                      //            dist6.rxd
		output wire        dist6_txd,                      //                 .txd
		input  wire        dist7_rxd,                      //            dist7.rxd
		output wire        dist7_txd,                      //                 .txd
		input  wire        dist8_rxd,                      //            dist8.rxd
		output wire        dist8_txd                       //                 .txd
	);

	wire         sys_pll_c0_clk;                                                                     // sys_pll:c0 -> [ACELEROMETRO_SPI:clk, ADC_DE0:clock, CPU:clk, CTRL_I2C:clk, DATA_IN_I2C:clk, DATA_OUT_I2C:clk, DIST1:clk, DIST2:clk, DIST3:clk, DIST4:clk, DIST5:clk, DIST6:clk, DIST7:clk, DIST8:clk, ENCODER_INT:clk, ENCODER_NORMAL:clk, EPCS:clk, FLAG_I2C:clk, GPS:clk, JTAG:clk, KEY:clk, LED:clk, MOTORES:clk, PWM1:clk, PWM2:clk, SDRAM:clk, SW:clk, XBEE:clk, irq_mapper:clk, mm_interconnect_0:sys_clk_clk_clk, rst_controller:clk, sys_id:clock, sys_timer:clk]
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;                                     // mm_interconnect_0:sys_id_control_slave_address -> sys_id:address
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;                                    // sys_id:readdata -> mm_interconnect_0:sys_id_control_slave_readdata
	wire  [15:0] mm_interconnect_0_dist4_s1_writedata;                                               // mm_interconnect_0:DIST4_s1_writedata -> DIST4:writedata
	wire   [2:0] mm_interconnect_0_dist4_s1_address;                                                 // mm_interconnect_0:DIST4_s1_address -> DIST4:address
	wire         mm_interconnect_0_dist4_s1_chipselect;                                              // mm_interconnect_0:DIST4_s1_chipselect -> DIST4:chipselect
	wire         mm_interconnect_0_dist4_s1_write;                                                   // mm_interconnect_0:DIST4_s1_write -> DIST4:write_n
	wire         mm_interconnect_0_dist4_s1_read;                                                    // mm_interconnect_0:DIST4_s1_read -> DIST4:read_n
	wire  [15:0] mm_interconnect_0_dist4_s1_readdata;                                                // DIST4:readdata -> mm_interconnect_0:DIST4_s1_readdata
	wire         mm_interconnect_0_dist4_s1_begintransfer;                                           // mm_interconnect_0:DIST4_s1_begintransfer -> DIST4:begintransfer
	wire  [15:0] mm_interconnect_0_dist7_s1_writedata;                                               // mm_interconnect_0:DIST7_s1_writedata -> DIST7:writedata
	wire   [2:0] mm_interconnect_0_dist7_s1_address;                                                 // mm_interconnect_0:DIST7_s1_address -> DIST7:address
	wire         mm_interconnect_0_dist7_s1_chipselect;                                              // mm_interconnect_0:DIST7_s1_chipselect -> DIST7:chipselect
	wire         mm_interconnect_0_dist7_s1_write;                                                   // mm_interconnect_0:DIST7_s1_write -> DIST7:write_n
	wire         mm_interconnect_0_dist7_s1_read;                                                    // mm_interconnect_0:DIST7_s1_read -> DIST7:read_n
	wire  [15:0] mm_interconnect_0_dist7_s1_readdata;                                                // DIST7:readdata -> mm_interconnect_0:DIST7_s1_readdata
	wire         mm_interconnect_0_dist7_s1_begintransfer;                                           // mm_interconnect_0:DIST7_s1_begintransfer -> DIST7:begintransfer
	wire  [31:0] mm_interconnect_0_encoder_int_s1_writedata;                                         // mm_interconnect_0:ENCODER_INT_s1_writedata -> ENCODER_INT:writedata
	wire   [1:0] mm_interconnect_0_encoder_int_s1_address;                                           // mm_interconnect_0:ENCODER_INT_s1_address -> ENCODER_INT:address
	wire         mm_interconnect_0_encoder_int_s1_chipselect;                                        // mm_interconnect_0:ENCODER_INT_s1_chipselect -> ENCODER_INT:chipselect
	wire         mm_interconnect_0_encoder_int_s1_write;                                             // mm_interconnect_0:ENCODER_INT_s1_write -> ENCODER_INT:write_n
	wire  [31:0] mm_interconnect_0_encoder_int_s1_readdata;                                          // ENCODER_INT:readdata -> mm_interconnect_0:ENCODER_INT_s1_readdata
	wire  [31:0] mm_interconnect_0_sys_pll_pll_slave_writedata;                                      // mm_interconnect_0:sys_pll_pll_slave_writedata -> sys_pll:writedata
	wire   [1:0] mm_interconnect_0_sys_pll_pll_slave_address;                                        // mm_interconnect_0:sys_pll_pll_slave_address -> sys_pll:address
	wire         mm_interconnect_0_sys_pll_pll_slave_write;                                          // mm_interconnect_0:sys_pll_pll_slave_write -> sys_pll:write
	wire         mm_interconnect_0_sys_pll_pll_slave_read;                                           // mm_interconnect_0:sys_pll_pll_slave_read -> sys_pll:read
	wire  [31:0] mm_interconnect_0_sys_pll_pll_slave_readdata;                                       // sys_pll:readdata -> mm_interconnect_0:sys_pll_pll_slave_readdata
	wire  [31:0] mm_interconnect_0_pwm1_s1_writedata;                                                // mm_interconnect_0:PWM1_s1_writedata -> PWM1:writedata
	wire   [1:0] mm_interconnect_0_pwm1_s1_address;                                                  // mm_interconnect_0:PWM1_s1_address -> PWM1:address
	wire         mm_interconnect_0_pwm1_s1_chipselect;                                               // mm_interconnect_0:PWM1_s1_chipselect -> PWM1:chipselect
	wire         mm_interconnect_0_pwm1_s1_write;                                                    // mm_interconnect_0:PWM1_s1_write -> PWM1:write_n
	wire  [31:0] mm_interconnect_0_pwm1_s1_readdata;                                                 // PWM1:readdata -> mm_interconnect_0:PWM1_s1_readdata
	wire   [1:0] mm_interconnect_0_flag_i2c_s1_address;                                              // mm_interconnect_0:FLAG_I2C_s1_address -> FLAG_I2C:address
	wire  [31:0] mm_interconnect_0_flag_i2c_s1_readdata;                                             // FLAG_I2C:readdata -> mm_interconnect_0:FLAG_I2C_s1_readdata
	wire   [1:0] mm_interconnect_0_encoder_normal_s1_address;                                        // mm_interconnect_0:ENCODER_NORMAL_s1_address -> ENCODER_NORMAL:address
	wire  [31:0] mm_interconnect_0_encoder_normal_s1_readdata;                                       // ENCODER_NORMAL:readdata -> mm_interconnect_0:ENCODER_NORMAL_s1_readdata
	wire  [15:0] mm_interconnect_0_dist5_s1_writedata;                                               // mm_interconnect_0:DIST5_s1_writedata -> DIST5:writedata
	wire   [2:0] mm_interconnect_0_dist5_s1_address;                                                 // mm_interconnect_0:DIST5_s1_address -> DIST5:address
	wire         mm_interconnect_0_dist5_s1_chipselect;                                              // mm_interconnect_0:DIST5_s1_chipselect -> DIST5:chipselect
	wire         mm_interconnect_0_dist5_s1_write;                                                   // mm_interconnect_0:DIST5_s1_write -> DIST5:write_n
	wire         mm_interconnect_0_dist5_s1_read;                                                    // mm_interconnect_0:DIST5_s1_read -> DIST5:read_n
	wire  [15:0] mm_interconnect_0_dist5_s1_readdata;                                                // DIST5:readdata -> mm_interconnect_0:DIST5_s1_readdata
	wire         mm_interconnect_0_dist5_s1_begintransfer;                                           // mm_interconnect_0:DIST5_s1_begintransfer -> DIST5:begintransfer
	wire  [15:0] mm_interconnect_0_xbee_s1_writedata;                                                // mm_interconnect_0:XBEE_s1_writedata -> XBEE:writedata
	wire   [2:0] mm_interconnect_0_xbee_s1_address;                                                  // mm_interconnect_0:XBEE_s1_address -> XBEE:address
	wire         mm_interconnect_0_xbee_s1_chipselect;                                               // mm_interconnect_0:XBEE_s1_chipselect -> XBEE:chipselect
	wire         mm_interconnect_0_xbee_s1_write;                                                    // mm_interconnect_0:XBEE_s1_write -> XBEE:write_n
	wire         mm_interconnect_0_xbee_s1_read;                                                     // mm_interconnect_0:XBEE_s1_read -> XBEE:read_n
	wire  [15:0] mm_interconnect_0_xbee_s1_readdata;                                                 // XBEE:readdata -> mm_interconnect_0:XBEE_s1_readdata
	wire         mm_interconnect_0_xbee_s1_begintransfer;                                            // mm_interconnect_0:XBEE_s1_begintransfer -> XBEE:begintransfer
	wire  [31:0] mm_interconnect_0_pwm2_s1_writedata;                                                // mm_interconnect_0:PWM2_s1_writedata -> PWM2:writedata
	wire   [1:0] mm_interconnect_0_pwm2_s1_address;                                                  // mm_interconnect_0:PWM2_s1_address -> PWM2:address
	wire         mm_interconnect_0_pwm2_s1_chipselect;                                               // mm_interconnect_0:PWM2_s1_chipselect -> PWM2:chipselect
	wire         mm_interconnect_0_pwm2_s1_write;                                                    // mm_interconnect_0:PWM2_s1_write -> PWM2:write_n
	wire  [31:0] mm_interconnect_0_pwm2_s1_readdata;                                                 // PWM2:readdata -> mm_interconnect_0:PWM2_s1_readdata
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_writedata;                                 // mm_interconnect_0:EPCS_epcs_control_port_writedata -> EPCS:writedata
	wire   [8:0] mm_interconnect_0_epcs_epcs_control_port_address;                                   // mm_interconnect_0:EPCS_epcs_control_port_address -> EPCS:address
	wire         mm_interconnect_0_epcs_epcs_control_port_chipselect;                                // mm_interconnect_0:EPCS_epcs_control_port_chipselect -> EPCS:chipselect
	wire         mm_interconnect_0_epcs_epcs_control_port_write;                                     // mm_interconnect_0:EPCS_epcs_control_port_write -> EPCS:write_n
	wire         mm_interconnect_0_epcs_epcs_control_port_read;                                      // mm_interconnect_0:EPCS_epcs_control_port_read -> EPCS:read_n
	wire  [31:0] mm_interconnect_0_epcs_epcs_control_port_readdata;                                  // EPCS:readdata -> mm_interconnect_0:EPCS_epcs_control_port_readdata
	wire   [1:0] mm_interconnect_0_data_in_i2c_s1_address;                                           // mm_interconnect_0:DATA_IN_I2C_s1_address -> DATA_IN_I2C:address
	wire  [31:0] mm_interconnect_0_data_in_i2c_s1_readdata;                                          // DATA_IN_I2C:readdata -> mm_interconnect_0:DATA_IN_I2C_s1_readdata
	wire  [31:0] mm_interconnect_0_led_s1_writedata;                                                 // mm_interconnect_0:LED_s1_writedata -> LED:writedata
	wire   [1:0] mm_interconnect_0_led_s1_address;                                                   // mm_interconnect_0:LED_s1_address -> LED:address
	wire         mm_interconnect_0_led_s1_chipselect;                                                // mm_interconnect_0:LED_s1_chipselect -> LED:chipselect
	wire         mm_interconnect_0_led_s1_write;                                                     // mm_interconnect_0:LED_s1_write -> LED:write_n
	wire  [31:0] mm_interconnect_0_led_s1_readdata;                                                  // LED:readdata -> mm_interconnect_0:LED_s1_readdata
	wire  [31:0] mm_interconnect_0_key_s1_writedata;                                                 // mm_interconnect_0:KEY_s1_writedata -> KEY:writedata
	wire   [1:0] mm_interconnect_0_key_s1_address;                                                   // mm_interconnect_0:KEY_s1_address -> KEY:address
	wire         mm_interconnect_0_key_s1_chipselect;                                                // mm_interconnect_0:KEY_s1_chipselect -> KEY:chipselect
	wire         mm_interconnect_0_key_s1_write;                                                     // mm_interconnect_0:KEY_s1_write -> KEY:write_n
	wire  [31:0] mm_interconnect_0_key_s1_readdata;                                                  // KEY:readdata -> mm_interconnect_0:KEY_s1_readdata
	wire  [15:0] mm_interconnect_0_dist2_s1_writedata;                                               // mm_interconnect_0:DIST2_s1_writedata -> DIST2:writedata
	wire   [2:0] mm_interconnect_0_dist2_s1_address;                                                 // mm_interconnect_0:DIST2_s1_address -> DIST2:address
	wire         mm_interconnect_0_dist2_s1_chipselect;                                              // mm_interconnect_0:DIST2_s1_chipselect -> DIST2:chipselect
	wire         mm_interconnect_0_dist2_s1_write;                                                   // mm_interconnect_0:DIST2_s1_write -> DIST2:write_n
	wire         mm_interconnect_0_dist2_s1_read;                                                    // mm_interconnect_0:DIST2_s1_read -> DIST2:read_n
	wire  [15:0] mm_interconnect_0_dist2_s1_readdata;                                                // DIST2:readdata -> mm_interconnect_0:DIST2_s1_readdata
	wire         mm_interconnect_0_dist2_s1_begintransfer;                                           // mm_interconnect_0:DIST2_s1_begintransfer -> DIST2:begintransfer
	wire  [15:0] mm_interconnect_0_dist1_s1_writedata;                                               // mm_interconnect_0:DIST1_s1_writedata -> DIST1:writedata
	wire   [2:0] mm_interconnect_0_dist1_s1_address;                                                 // mm_interconnect_0:DIST1_s1_address -> DIST1:address
	wire         mm_interconnect_0_dist1_s1_chipselect;                                              // mm_interconnect_0:DIST1_s1_chipselect -> DIST1:chipselect
	wire         mm_interconnect_0_dist1_s1_write;                                                   // mm_interconnect_0:DIST1_s1_write -> DIST1:write_n
	wire         mm_interconnect_0_dist1_s1_read;                                                    // mm_interconnect_0:DIST1_s1_read -> DIST1:read_n
	wire  [15:0] mm_interconnect_0_dist1_s1_readdata;                                                // DIST1:readdata -> mm_interconnect_0:DIST1_s1_readdata
	wire         mm_interconnect_0_dist1_s1_begintransfer;                                           // mm_interconnect_0:DIST1_s1_begintransfer -> DIST1:begintransfer
	wire  [15:0] mm_interconnect_0_dist8_s1_writedata;                                               // mm_interconnect_0:DIST8_s1_writedata -> DIST8:writedata
	wire   [2:0] mm_interconnect_0_dist8_s1_address;                                                 // mm_interconnect_0:DIST8_s1_address -> DIST8:address
	wire         mm_interconnect_0_dist8_s1_chipselect;                                              // mm_interconnect_0:DIST8_s1_chipselect -> DIST8:chipselect
	wire         mm_interconnect_0_dist8_s1_write;                                                   // mm_interconnect_0:DIST8_s1_write -> DIST8:write_n
	wire         mm_interconnect_0_dist8_s1_read;                                                    // mm_interconnect_0:DIST8_s1_read -> DIST8:read_n
	wire  [15:0] mm_interconnect_0_dist8_s1_readdata;                                                // DIST8:readdata -> mm_interconnect_0:DIST8_s1_readdata
	wire         mm_interconnect_0_dist8_s1_begintransfer;                                           // mm_interconnect_0:DIST8_s1_begintransfer -> DIST8:begintransfer
	wire  [15:0] mm_interconnect_0_gps_s1_writedata;                                                 // mm_interconnect_0:GPS_s1_writedata -> GPS:writedata
	wire   [2:0] mm_interconnect_0_gps_s1_address;                                                   // mm_interconnect_0:GPS_s1_address -> GPS:address
	wire         mm_interconnect_0_gps_s1_chipselect;                                                // mm_interconnect_0:GPS_s1_chipselect -> GPS:chipselect
	wire         mm_interconnect_0_gps_s1_write;                                                     // mm_interconnect_0:GPS_s1_write -> GPS:write_n
	wire         mm_interconnect_0_gps_s1_read;                                                      // mm_interconnect_0:GPS_s1_read -> GPS:read_n
	wire  [15:0] mm_interconnect_0_gps_s1_readdata;                                                  // GPS:readdata -> mm_interconnect_0:GPS_s1_readdata
	wire         mm_interconnect_0_gps_s1_begintransfer;                                             // mm_interconnect_0:GPS_s1_begintransfer -> GPS:begintransfer
	wire  [15:0] mm_interconnect_0_sys_timer_s1_writedata;                                           // mm_interconnect_0:sys_timer_s1_writedata -> sys_timer:writedata
	wire   [2:0] mm_interconnect_0_sys_timer_s1_address;                                             // mm_interconnect_0:sys_timer_s1_address -> sys_timer:address
	wire         mm_interconnect_0_sys_timer_s1_chipselect;                                          // mm_interconnect_0:sys_timer_s1_chipselect -> sys_timer:chipselect
	wire         mm_interconnect_0_sys_timer_s1_write;                                               // mm_interconnect_0:sys_timer_s1_write -> sys_timer:write_n
	wire  [15:0] mm_interconnect_0_sys_timer_s1_readdata;                                            // sys_timer:readdata -> mm_interconnect_0:sys_timer_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                                             // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [15:0] mm_interconnect_0_sdram_s1_writedata;                                               // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire  [23:0] mm_interconnect_0_sdram_s1_address;                                                 // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_chipselect;                                              // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire         mm_interconnect_0_sdram_s1_write;                                                   // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire         mm_interconnect_0_sdram_s1_read;                                                    // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire  [15:0] mm_interconnect_0_sdram_s1_readdata;                                                // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                                           // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire   [1:0] mm_interconnect_0_sdram_s1_byteenable;                                              // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_cpu_jtag_debug_module_waitrequest;                                // CPU:jtag_debug_module_waitrequest -> mm_interconnect_0:CPU_jtag_debug_module_waitrequest
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;                                  // mm_interconnect_0:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	wire   [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;                                    // mm_interconnect_0:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	wire         mm_interconnect_0_cpu_jtag_debug_module_write;                                      // mm_interconnect_0:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	wire         mm_interconnect_0_cpu_jtag_debug_module_read;                                       // mm_interconnect_0:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	wire  [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;                                   // CPU:jtag_debug_module_readdata -> mm_interconnect_0:CPU_jtag_debug_module_readdata
	wire         mm_interconnect_0_cpu_jtag_debug_module_debugaccess;                                // mm_interconnect_0:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	wire   [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;                                 // mm_interconnect_0:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	wire  [15:0] mm_interconnect_0_dist3_s1_writedata;                                               // mm_interconnect_0:DIST3_s1_writedata -> DIST3:writedata
	wire   [2:0] mm_interconnect_0_dist3_s1_address;                                                 // mm_interconnect_0:DIST3_s1_address -> DIST3:address
	wire         mm_interconnect_0_dist3_s1_chipselect;                                              // mm_interconnect_0:DIST3_s1_chipselect -> DIST3:chipselect
	wire         mm_interconnect_0_dist3_s1_write;                                                   // mm_interconnect_0:DIST3_s1_write -> DIST3:write_n
	wire         mm_interconnect_0_dist3_s1_read;                                                    // mm_interconnect_0:DIST3_s1_read -> DIST3:read_n
	wire  [15:0] mm_interconnect_0_dist3_s1_readdata;                                                // DIST3:readdata -> mm_interconnect_0:DIST3_s1_readdata
	wire         mm_interconnect_0_dist3_s1_begintransfer;                                           // mm_interconnect_0:DIST3_s1_begintransfer -> DIST3:begintransfer
	wire         cpu_instruction_master_waitrequest;                                                 // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [26:0] cpu_instruction_master_address;                                                     // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                                                        // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire  [31:0] cpu_instruction_master_readdata;                                                    // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_readdatavalid;                                               // mm_interconnect_0:CPU_instruction_master_readdatavalid -> CPU:i_readdatavalid
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest;                               // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;                                 // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;                                   // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;                                // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;                                     // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;                                      // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;                                  // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         cpu_data_master_waitrequest;                                                        // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire  [31:0] cpu_data_master_writedata;                                                          // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [26:0] cpu_data_master_address;                                                            // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire         cpu_data_master_write;                                                              // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire         cpu_data_master_read;                                                               // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire  [31:0] cpu_data_master_readdata;                                                           // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_debugaccess;                                                        // CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire   [3:0] cpu_data_master_byteenable;                                                         // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_waitrequest; // ACELEROMETRO_SPI:waitrequest -> mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_waitrequest
	wire   [7:0] mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_writedata;   // mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_writedata -> ACELEROMETRO_SPI:writedata
	wire   [0:0] mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_address;     // mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_address -> ACELEROMETRO_SPI:address
	wire         mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_write;       // mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_write -> ACELEROMETRO_SPI:write
	wire         mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_read;        // mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_read -> ACELEROMETRO_SPI:read
	wire   [7:0] mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_readdata;    // ACELEROMETRO_SPI:readdata -> mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_readdata
	wire   [0:0] mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_byteenable;  // mm_interconnect_0:ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_byteenable -> ACELEROMETRO_SPI:byteenable
	wire  [15:0] mm_interconnect_0_dist6_s1_writedata;                                               // mm_interconnect_0:DIST6_s1_writedata -> DIST6:writedata
	wire   [2:0] mm_interconnect_0_dist6_s1_address;                                                 // mm_interconnect_0:DIST6_s1_address -> DIST6:address
	wire         mm_interconnect_0_dist6_s1_chipselect;                                              // mm_interconnect_0:DIST6_s1_chipselect -> DIST6:chipselect
	wire         mm_interconnect_0_dist6_s1_write;                                                   // mm_interconnect_0:DIST6_s1_write -> DIST6:write_n
	wire         mm_interconnect_0_dist6_s1_read;                                                    // mm_interconnect_0:DIST6_s1_read -> DIST6:read_n
	wire  [15:0] mm_interconnect_0_dist6_s1_readdata;                                                // DIST6:readdata -> mm_interconnect_0:DIST6_s1_readdata
	wire         mm_interconnect_0_dist6_s1_begintransfer;                                           // mm_interconnect_0:DIST6_s1_begintransfer -> DIST6:begintransfer
	wire  [31:0] mm_interconnect_0_motores_s1_writedata;                                             // mm_interconnect_0:MOTORES_s1_writedata -> MOTORES:writedata
	wire   [1:0] mm_interconnect_0_motores_s1_address;                                               // mm_interconnect_0:MOTORES_s1_address -> MOTORES:address
	wire         mm_interconnect_0_motores_s1_chipselect;                                            // mm_interconnect_0:MOTORES_s1_chipselect -> MOTORES:chipselect
	wire         mm_interconnect_0_motores_s1_write;                                                 // mm_interconnect_0:MOTORES_s1_write -> MOTORES:write_n
	wire  [31:0] mm_interconnect_0_motores_s1_readdata;                                              // MOTORES:readdata -> mm_interconnect_0:MOTORES_s1_readdata
	wire   [1:0] mm_interconnect_0_sw_s1_address;                                                    // mm_interconnect_0:SW_s1_address -> SW:address
	wire  [31:0] mm_interconnect_0_sw_s1_readdata;                                                   // SW:readdata -> mm_interconnect_0:SW_s1_readdata
	wire         mm_interconnect_0_adc_de0_adc_slave_waitrequest;                                    // ADC_DE0:waitrequest -> mm_interconnect_0:ADC_DE0_adc_slave_waitrequest
	wire  [31:0] mm_interconnect_0_adc_de0_adc_slave_writedata;                                      // mm_interconnect_0:ADC_DE0_adc_slave_writedata -> ADC_DE0:writedata
	wire   [2:0] mm_interconnect_0_adc_de0_adc_slave_address;                                        // mm_interconnect_0:ADC_DE0_adc_slave_address -> ADC_DE0:address
	wire         mm_interconnect_0_adc_de0_adc_slave_write;                                          // mm_interconnect_0:ADC_DE0_adc_slave_write -> ADC_DE0:write
	wire         mm_interconnect_0_adc_de0_adc_slave_read;                                           // mm_interconnect_0:ADC_DE0_adc_slave_read -> ADC_DE0:read
	wire  [31:0] mm_interconnect_0_adc_de0_adc_slave_readdata;                                       // ADC_DE0:readdata -> mm_interconnect_0:ADC_DE0_adc_slave_readdata
	wire  [31:0] mm_interconnect_0_data_out_i2c_s1_writedata;                                        // mm_interconnect_0:DATA_OUT_I2C_s1_writedata -> DATA_OUT_I2C:writedata
	wire   [1:0] mm_interconnect_0_data_out_i2c_s1_address;                                          // mm_interconnect_0:DATA_OUT_I2C_s1_address -> DATA_OUT_I2C:address
	wire         mm_interconnect_0_data_out_i2c_s1_chipselect;                                       // mm_interconnect_0:DATA_OUT_I2C_s1_chipselect -> DATA_OUT_I2C:chipselect
	wire         mm_interconnect_0_data_out_i2c_s1_write;                                            // mm_interconnect_0:DATA_OUT_I2C_s1_write -> DATA_OUT_I2C:write_n
	wire  [31:0] mm_interconnect_0_data_out_i2c_s1_readdata;                                         // DATA_OUT_I2C:readdata -> mm_interconnect_0:DATA_OUT_I2C_s1_readdata
	wire  [31:0] mm_interconnect_0_ctrl_i2c_s1_writedata;                                            // mm_interconnect_0:CTRL_I2C_s1_writedata -> CTRL_I2C:writedata
	wire   [1:0] mm_interconnect_0_ctrl_i2c_s1_address;                                              // mm_interconnect_0:CTRL_I2C_s1_address -> CTRL_I2C:address
	wire         mm_interconnect_0_ctrl_i2c_s1_chipselect;                                           // mm_interconnect_0:CTRL_I2C_s1_chipselect -> CTRL_I2C:chipselect
	wire         mm_interconnect_0_ctrl_i2c_s1_write;                                                // mm_interconnect_0:CTRL_I2C_s1_write -> CTRL_I2C:write_n
	wire  [31:0] mm_interconnect_0_ctrl_i2c_s1_readdata;                                             // CTRL_I2C:readdata -> mm_interconnect_0:CTRL_I2C_s1_readdata
	wire         irq_mapper_receiver0_irq;                                                           // EPCS:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                                           // sys_timer:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                                                           // JTAG:av_irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                                                           // KEY:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                                                           // ENCODER_INT:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                                                           // ACELEROMETRO_SPI:irq -> irq_mapper:receiver5_irq
	wire         irq_mapper_receiver6_irq;                                                           // GPS:irq -> irq_mapper:receiver6_irq
	wire         irq_mapper_receiver7_irq;                                                           // XBEE:irq -> irq_mapper:receiver7_irq
	wire         irq_mapper_receiver8_irq;                                                           // DIST1:irq -> irq_mapper:receiver8_irq
	wire         irq_mapper_receiver9_irq;                                                           // DIST2:irq -> irq_mapper:receiver9_irq
	wire         irq_mapper_receiver10_irq;                                                          // DIST3:irq -> irq_mapper:receiver10_irq
	wire         irq_mapper_receiver11_irq;                                                          // DIST4:irq -> irq_mapper:receiver11_irq
	wire         irq_mapper_receiver12_irq;                                                          // DIST5:irq -> irq_mapper:receiver12_irq
	wire         irq_mapper_receiver13_irq;                                                          // DIST6:irq -> irq_mapper:receiver13_irq
	wire         irq_mapper_receiver14_irq;                                                          // DIST7:irq -> irq_mapper:receiver14_irq
	wire         irq_mapper_receiver15_irq;                                                          // DIST8:irq -> irq_mapper:receiver15_irq
	wire  [31:0] cpu_d_irq_irq;                                                                      // irq_mapper:sender_irq -> CPU:d_irq
	wire         rst_controller_reset_out_reset;                                                     // rst_controller:reset_out -> [ACELEROMETRO_SPI:reset, ADC_DE0:reset, CPU:reset_n, CTRL_I2C:reset_n, DATA_IN_I2C:reset_n, DATA_OUT_I2C:reset_n, DIST1:reset_n, DIST2:reset_n, DIST3:reset_n, DIST4:reset_n, DIST5:reset_n, DIST6:reset_n, DIST7:reset_n, DIST8:reset_n, ENCODER_INT:reset_n, ENCODER_NORMAL:reset_n, EPCS:reset_n, FLAG_I2C:reset_n, GPS:reset_n, JTAG:rst_n, KEY:reset_n, LED:reset_n, MOTORES:reset_n, PWM1:reset_n, PWM2:reset_n, SDRAM:reset_n, SW:reset_n, XBEE:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_n_reset_bridge_in_reset_reset, rst_translator:in_reset, sys_id:reset_n, sys_timer:reset_n]
	wire         rst_controller_reset_out_reset_req;                                                 // rst_controller:reset_req -> [CPU:reset_req, EPCS:reset_req, rst_translator:reset_req_in]
	wire         cpu_jtag_debug_module_reset_reset;                                                  // CPU:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1, rst_controller_002:reset_in1, rst_controller_003:reset_in1]
	wire         rst_controller_001_reset_out_reset;                                                 // rst_controller_001:reset_out -> [mm_interconnect_0:sys_pll_inclk_interface_reset_reset_bridge_in_reset_reset, sys_pll:reset]
	wire         rst_controller_002_reset_out_reset;                                                 // rst_controller_002:reset_out -> [rst_controller:reset_in2, rst_controller_001:reset_in2]
	wire         rst_controller_003_reset_out_reset;                                                 // rst_controller_003:reset_out -> [rst_controller:reset_in3, rst_controller_001:reset_in3]

	NIOS_CPU cpu (
		.clk                                   (sys_pll_c0_clk),                                      //                       clk.clk
		.reset_n                               (~rst_controller_reset_out_reset),                     //                   reset_n.reset_n
		.reset_req                             (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	NIOS_sys_id sys_id (
		.clock    (sys_pll_c0_clk),                                  //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	NIOS_SDRAM sdram (
		.clk            (sys_pll_c0_clk),                           //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_addr),                               //  wire.export
		.zs_ba          (sdram_ba),                                 //      .export
		.zs_cas_n       (sdram_cas_n),                              //      .export
		.zs_cke         (sdram_cke),                                //      .export
		.zs_cs_n        (sdram_cs_n),                               //      .export
		.zs_dq          (sdram_dq),                                 //      .export
		.zs_dqm         (sdram_dqm),                                //      .export
		.zs_ras_n       (sdram_ras_n),                              //      .export
		.zs_we_n        (sdram_we_n)                                //      .export
	);

	NIOS_EPCS epcs (
		.clk           (sys_pll_c0_clk),                                      //               clk.clk
		.reset_n       (~rst_controller_reset_out_reset),                     //             reset.reset_n
		.reset_req     (rst_controller_reset_out_reset_req),                  //                  .reset_req
		.address       (mm_interconnect_0_epcs_epcs_control_port_address),    // epcs_control_port.address
		.chipselect    (mm_interconnect_0_epcs_epcs_control_port_chipselect), //                  .chipselect
		.dataavailable (),                                                    //                  .dataavailable
		.endofpacket   (),                                                    //                  .endofpacket
		.read_n        (~mm_interconnect_0_epcs_epcs_control_port_read),      //                  .read_n
		.readdata      (mm_interconnect_0_epcs_epcs_control_port_readdata),   //                  .readdata
		.readyfordata  (),                                                    //                  .readyfordata
		.write_n       (~mm_interconnect_0_epcs_epcs_control_port_write),     //                  .write_n
		.writedata     (mm_interconnect_0_epcs_epcs_control_port_writedata),  //                  .writedata
		.irq           (irq_mapper_receiver0_irq),                            //               irq.irq
		.dclk          (epcs_dclk),                                           //          external.export
		.sce           (epcs_sce),                                            //                  .export
		.sdo           (epcs_sdo),                                            //                  .export
		.data0         (epcs_data0)                                           //                  .export
	);

	NIOS_sys_timer sys_timer (
		.clk        (sys_pll_c0_clk),                            //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_sys_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_sys_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_sys_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_sys_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_sys_timer_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                   //   irq.irq
	);

	NIOS_LED led (
		.clk        (sys_pll_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_led_s1_readdata),   //                    .readdata
		.out_port   (led_export)                           // external_connection.export
	);

	NIOS_SW sw (
		.clk      (sys_pll_c0_clk),                   //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),  //               reset.reset_n
		.address  (mm_interconnect_0_sw_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_sw_s1_readdata), //                    .readdata
		.in_port  (sw_export)                         // external_connection.export
	);

	NIOS_KEY key (
		.clk        (sys_pll_c0_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_0_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_key_s1_readdata),   //                    .readdata
		.in_port    (key_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)             //                 irq.irq
	);

	NIOS_JTAG jtag (
		.clk            (sys_pll_c0_clk),                                       //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver2_irq)                              //               irq.irq
	);

	NIOS_sys_pll sys_pll (
		.clk       (clk_clk),                                       //       inclk_interface.clk
		.reset     (rst_controller_001_reset_out_reset),            // inclk_interface_reset.reset
		.read      (mm_interconnect_0_sys_pll_pll_slave_read),      //             pll_slave.read
		.write     (mm_interconnect_0_sys_pll_pll_slave_write),     //                      .write
		.address   (mm_interconnect_0_sys_pll_pll_slave_address),   //                      .address
		.readdata  (mm_interconnect_0_sys_pll_pll_slave_readdata),  //                      .readdata
		.writedata (mm_interconnect_0_sys_pll_pll_slave_writedata), //                      .writedata
		.c0        (sys_pll_c0_clk),                                //                    c0.clk
		.c1        (ram_clk_clk),                                   //                    c1.clk
		.areset    (),                                              //        areset_conduit.export
		.locked    (),                                              //        locked_conduit.export
		.phasedone ()                                               //     phasedone_conduit.export
	);

	NIOS_ACELEROMETRO_SPI acelerometro_spi (
		.clk           (sys_pll_c0_clk),                                                                     //                         clock_reset.clk
		.reset         (rst_controller_reset_out_reset),                                                     //                   clock_reset_reset.reset
		.address       (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_address),     // avalon_accelerometer_spi_mode_slave.address
		.byteenable    (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_byteenable),  //                                    .byteenable
		.read          (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_read),        //                                    .read
		.write         (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_write),       //                                    .write
		.writedata     (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_writedata),   //                                    .writedata
		.readdata      (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_readdata),    //                                    .readdata
		.waitrequest   (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_waitrequest), //                                    .waitrequest
		.irq           (irq_mapper_receiver5_irq),                                                           //                           interrupt.irq
		.I2C_SDAT      (acelerometro_spi_I2C_SDAT),                                                          //                  external_interface.export
		.I2C_SCLK      (acelerometro_spi_I2C_SCLK),                                                          //                                    .export
		.G_SENSOR_CS_N (acelerometro_spi_G_SENSOR_CS_N),                                                     //                                    .export
		.G_SENSOR_INT  (acelerometro_spi_G_SENSOR_INT)                                                       //                                    .export
	);

	NIOS_ADC_DE0 adc_de0 (
		.clock       (sys_pll_c0_clk),                                  //                clk.clk
		.reset       (rst_controller_reset_out_reset),                  //              reset.reset
		.write       (mm_interconnect_0_adc_de0_adc_slave_write),       //          adc_slave.write
		.readdata    (mm_interconnect_0_adc_de0_adc_slave_readdata),    //                   .readdata
		.writedata   (mm_interconnect_0_adc_de0_adc_slave_writedata),   //                   .writedata
		.address     (mm_interconnect_0_adc_de0_adc_slave_address),     //                   .address
		.waitrequest (mm_interconnect_0_adc_de0_adc_slave_waitrequest), //                   .waitrequest
		.read        (mm_interconnect_0_adc_de0_adc_slave_read),        //                   .read
		.adc_sclk    (adc_sclk),                                        // external_interface.export
		.adc_cs_n    (adc_cs_n),                                        //                   .export
		.adc_dout    (adc_dout),                                        //                   .export
		.adc_din     (adc_din)                                          //                   .export
	);

	NIOS_ENCODER_INT encoder_int (
		.clk        (sys_pll_c0_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_encoder_int_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_encoder_int_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_encoder_int_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_encoder_int_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_encoder_int_s1_readdata),   //                    .readdata
		.in_port    (encoder_int_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                     //                 irq.irq
	);

	NIOS_SW encoder_normal (
		.clk      (sys_pll_c0_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address  (mm_interconnect_0_encoder_normal_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_encoder_normal_s1_readdata), //                    .readdata
		.in_port  (encoder_normal_export)                         // external_connection.export
	);

	NIOS_MOTORES motores (
		.clk        (sys_pll_c0_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_motores_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_motores_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_motores_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_motores_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_motores_s1_readdata),   //                    .readdata
		.out_port   (motores_export)                           // external_connection.export
	);

	NIOS_LED pwm1 (
		.clk        (sys_pll_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_pwm1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pwm1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pwm1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pwm1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pwm1_s1_readdata),   //                    .readdata
		.out_port   (pwm1_export)                           // external_connection.export
	);

	NIOS_LED pwm2 (
		.clk        (sys_pll_c0_clk),                       //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_pwm2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_pwm2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_pwm2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_pwm2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_pwm2_s1_readdata),   //                    .readdata
		.out_port   (pwm2_export)                           // external_connection.export
	);

	NIOS_CTRL_I2C ctrl_i2c (
		.clk        (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_ctrl_i2c_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ctrl_i2c_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ctrl_i2c_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ctrl_i2c_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ctrl_i2c_s1_readdata),   //                    .readdata
		.out_port   (ctrl_i2c_export)                           // external_connection.export
	);

	NIOS_LED data_out_i2c (
		.clk        (sys_pll_c0_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),              //               reset.reset_n
		.address    (mm_interconnect_0_data_out_i2c_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_data_out_i2c_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_data_out_i2c_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_data_out_i2c_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_data_out_i2c_s1_readdata),   //                    .readdata
		.out_port   (data_out_i2c_export)                           // external_connection.export
	);

	NIOS_DATA_IN_I2C data_in_i2c (
		.clk      (sys_pll_c0_clk),                            //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),           //               reset.reset_n
		.address  (mm_interconnect_0_data_in_i2c_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_data_in_i2c_s1_readdata), //                    .readdata
		.in_port  (data_in_i2c_export)                         // external_connection.export
	);

	NIOS_FLAG_I2C flag_i2c (
		.clk      (sys_pll_c0_clk),                         //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_flag_i2c_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_flag_i2c_s1_readdata), //                    .readdata
		.in_port  (flag_i2c_export)                         // external_connection.export
	);

	NIOS_GPS gps (
		.clk           (sys_pll_c0_clk),                         //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address       (mm_interconnect_0_gps_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_gps_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_gps_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_gps_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_gps_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_gps_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_gps_s1_readdata),      //                    .readdata
		.dataavailable (),                                       //                    .dataavailable
		.readyfordata  (),                                       //                    .readyfordata
		.rxd           (gps_rxd),                                // external_connection.export
		.txd           (gps_txd),                                //                    .export
		.irq           (irq_mapper_receiver6_irq)                //                 irq.irq
	);

	NIOS_GPS xbee (
		.clk           (sys_pll_c0_clk),                          //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_xbee_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_xbee_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_xbee_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_xbee_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_xbee_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_xbee_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_xbee_s1_readdata),      //                    .readdata
		.dataavailable (),                                        //                    .dataavailable
		.readyfordata  (),                                        //                    .readyfordata
		.rxd           (xbee_rxd),                                // external_connection.export
		.txd           (xbee_txd),                                //                    .export
		.irq           (irq_mapper_receiver7_irq)                 //                 irq.irq
	);

	NIOS_GPS dist1 (
		.clk           (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_dist1_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_dist1_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_dist1_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_dist1_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_dist1_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_dist1_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_dist1_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (dist1_rxd),                                // external_connection.export
		.txd           (dist1_txd),                                //                    .export
		.irq           (irq_mapper_receiver8_irq)                  //                 irq.irq
	);

	NIOS_GPS dist2 (
		.clk           (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_dist2_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_dist2_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_dist2_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_dist2_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_dist2_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_dist2_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_dist2_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (dist2_rxd),                                // external_connection.export
		.txd           (dist2_txd),                                //                    .export
		.irq           (irq_mapper_receiver9_irq)                  //                 irq.irq
	);

	NIOS_GPS dist3 (
		.clk           (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_dist3_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_dist3_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_dist3_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_dist3_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_dist3_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_dist3_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_dist3_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (dist3_rxd),                                // external_connection.export
		.txd           (dist3_txd),                                //                    .export
		.irq           (irq_mapper_receiver10_irq)                 //                 irq.irq
	);

	NIOS_GPS dist4 (
		.clk           (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_dist4_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_dist4_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_dist4_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_dist4_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_dist4_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_dist4_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_dist4_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (dist4_rxd),                                // external_connection.export
		.txd           (dist4_txd),                                //                    .export
		.irq           (irq_mapper_receiver11_irq)                 //                 irq.irq
	);

	NIOS_GPS dist5 (
		.clk           (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_dist5_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_dist5_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_dist5_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_dist5_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_dist5_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_dist5_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_dist5_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (dist5_rxd),                                // external_connection.export
		.txd           (dist5_txd),                                //                    .export
		.irq           (irq_mapper_receiver12_irq)                 //                 irq.irq
	);

	NIOS_GPS dist6 (
		.clk           (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_dist6_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_dist6_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_dist6_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_dist6_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_dist6_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_dist6_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_dist6_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (dist6_rxd),                                // external_connection.export
		.txd           (dist6_txd),                                //                    .export
		.irq           (irq_mapper_receiver13_irq)                 //                 irq.irq
	);

	NIOS_GPS dist7 (
		.clk           (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_dist7_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_dist7_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_dist7_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_dist7_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_dist7_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_dist7_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_dist7_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (dist7_rxd),                                // external_connection.export
		.txd           (dist7_txd),                                //                    .export
		.irq           (irq_mapper_receiver14_irq)                 //                 irq.irq
	);

	NIOS_GPS dist8 (
		.clk           (sys_pll_c0_clk),                           //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),          //               reset.reset_n
		.address       (mm_interconnect_0_dist8_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_dist8_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_dist8_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_dist8_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_dist8_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_dist8_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_dist8_s1_readdata),      //                    .readdata
		.dataavailable (),                                         //                    .dataavailable
		.readyfordata  (),                                         //                    .readyfordata
		.rxd           (dist8_rxd),                                // external_connection.export
		.txd           (dist8_txd),                                //                    .export
		.irq           (irq_mapper_receiver15_irq)                 //                 irq.irq
	);

	NIOS_mm_interconnect_0 mm_interconnect_0 (
		.clk_50_clk_clk                                                   (clk_clk),                                                                            //                                           clk_50_clk.clk
		.sys_clk_clk_clk                                                  (sys_pll_c0_clk),                                                                     //                                          sys_clk_clk.clk
		.CPU_reset_n_reset_bridge_in_reset_reset                          (rst_controller_reset_out_reset),                                                     //                    CPU_reset_n_reset_bridge_in_reset.reset
		.sys_pll_inclk_interface_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                                                 //  sys_pll_inclk_interface_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                                          (cpu_data_master_address),                                                            //                                      CPU_data_master.address
		.CPU_data_master_waitrequest                                      (cpu_data_master_waitrequest),                                                        //                                                     .waitrequest
		.CPU_data_master_byteenable                                       (cpu_data_master_byteenable),                                                         //                                                     .byteenable
		.CPU_data_master_read                                             (cpu_data_master_read),                                                               //                                                     .read
		.CPU_data_master_readdata                                         (cpu_data_master_readdata),                                                           //                                                     .readdata
		.CPU_data_master_write                                            (cpu_data_master_write),                                                              //                                                     .write
		.CPU_data_master_writedata                                        (cpu_data_master_writedata),                                                          //                                                     .writedata
		.CPU_data_master_debugaccess                                      (cpu_data_master_debugaccess),                                                        //                                                     .debugaccess
		.CPU_instruction_master_address                                   (cpu_instruction_master_address),                                                     //                               CPU_instruction_master.address
		.CPU_instruction_master_waitrequest                               (cpu_instruction_master_waitrequest),                                                 //                                                     .waitrequest
		.CPU_instruction_master_read                                      (cpu_instruction_master_read),                                                        //                                                     .read
		.CPU_instruction_master_readdata                                  (cpu_instruction_master_readdata),                                                    //                                                     .readdata
		.CPU_instruction_master_readdatavalid                             (cpu_instruction_master_readdatavalid),                                               //                                                     .readdatavalid
		.ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_address     (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_address),     // ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave.address
		.ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_write       (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_write),       //                                                     .write
		.ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_read        (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_read),        //                                                     .read
		.ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_readdata    (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_readdata),    //                                                     .readdata
		.ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_writedata   (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_writedata),   //                                                     .writedata
		.ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_byteenable  (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_byteenable),  //                                                     .byteenable
		.ACELEROMETRO_SPI_avalon_accelerometer_spi_mode_slave_waitrequest (mm_interconnect_0_acelerometro_spi_avalon_accelerometer_spi_mode_slave_waitrequest), //                                                     .waitrequest
		.ADC_DE0_adc_slave_address                                        (mm_interconnect_0_adc_de0_adc_slave_address),                                        //                                    ADC_DE0_adc_slave.address
		.ADC_DE0_adc_slave_write                                          (mm_interconnect_0_adc_de0_adc_slave_write),                                          //                                                     .write
		.ADC_DE0_adc_slave_read                                           (mm_interconnect_0_adc_de0_adc_slave_read),                                           //                                                     .read
		.ADC_DE0_adc_slave_readdata                                       (mm_interconnect_0_adc_de0_adc_slave_readdata),                                       //                                                     .readdata
		.ADC_DE0_adc_slave_writedata                                      (mm_interconnect_0_adc_de0_adc_slave_writedata),                                      //                                                     .writedata
		.ADC_DE0_adc_slave_waitrequest                                    (mm_interconnect_0_adc_de0_adc_slave_waitrequest),                                    //                                                     .waitrequest
		.CPU_jtag_debug_module_address                                    (mm_interconnect_0_cpu_jtag_debug_module_address),                                    //                                CPU_jtag_debug_module.address
		.CPU_jtag_debug_module_write                                      (mm_interconnect_0_cpu_jtag_debug_module_write),                                      //                                                     .write
		.CPU_jtag_debug_module_read                                       (mm_interconnect_0_cpu_jtag_debug_module_read),                                       //                                                     .read
		.CPU_jtag_debug_module_readdata                                   (mm_interconnect_0_cpu_jtag_debug_module_readdata),                                   //                                                     .readdata
		.CPU_jtag_debug_module_writedata                                  (mm_interconnect_0_cpu_jtag_debug_module_writedata),                                  //                                                     .writedata
		.CPU_jtag_debug_module_byteenable                                 (mm_interconnect_0_cpu_jtag_debug_module_byteenable),                                 //                                                     .byteenable
		.CPU_jtag_debug_module_waitrequest                                (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),                                //                                                     .waitrequest
		.CPU_jtag_debug_module_debugaccess                                (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),                                //                                                     .debugaccess
		.CTRL_I2C_s1_address                                              (mm_interconnect_0_ctrl_i2c_s1_address),                                              //                                          CTRL_I2C_s1.address
		.CTRL_I2C_s1_write                                                (mm_interconnect_0_ctrl_i2c_s1_write),                                                //                                                     .write
		.CTRL_I2C_s1_readdata                                             (mm_interconnect_0_ctrl_i2c_s1_readdata),                                             //                                                     .readdata
		.CTRL_I2C_s1_writedata                                            (mm_interconnect_0_ctrl_i2c_s1_writedata),                                            //                                                     .writedata
		.CTRL_I2C_s1_chipselect                                           (mm_interconnect_0_ctrl_i2c_s1_chipselect),                                           //                                                     .chipselect
		.DATA_IN_I2C_s1_address                                           (mm_interconnect_0_data_in_i2c_s1_address),                                           //                                       DATA_IN_I2C_s1.address
		.DATA_IN_I2C_s1_readdata                                          (mm_interconnect_0_data_in_i2c_s1_readdata),                                          //                                                     .readdata
		.DATA_OUT_I2C_s1_address                                          (mm_interconnect_0_data_out_i2c_s1_address),                                          //                                      DATA_OUT_I2C_s1.address
		.DATA_OUT_I2C_s1_write                                            (mm_interconnect_0_data_out_i2c_s1_write),                                            //                                                     .write
		.DATA_OUT_I2C_s1_readdata                                         (mm_interconnect_0_data_out_i2c_s1_readdata),                                         //                                                     .readdata
		.DATA_OUT_I2C_s1_writedata                                        (mm_interconnect_0_data_out_i2c_s1_writedata),                                        //                                                     .writedata
		.DATA_OUT_I2C_s1_chipselect                                       (mm_interconnect_0_data_out_i2c_s1_chipselect),                                       //                                                     .chipselect
		.DIST1_s1_address                                                 (mm_interconnect_0_dist1_s1_address),                                                 //                                             DIST1_s1.address
		.DIST1_s1_write                                                   (mm_interconnect_0_dist1_s1_write),                                                   //                                                     .write
		.DIST1_s1_read                                                    (mm_interconnect_0_dist1_s1_read),                                                    //                                                     .read
		.DIST1_s1_readdata                                                (mm_interconnect_0_dist1_s1_readdata),                                                //                                                     .readdata
		.DIST1_s1_writedata                                               (mm_interconnect_0_dist1_s1_writedata),                                               //                                                     .writedata
		.DIST1_s1_begintransfer                                           (mm_interconnect_0_dist1_s1_begintransfer),                                           //                                                     .begintransfer
		.DIST1_s1_chipselect                                              (mm_interconnect_0_dist1_s1_chipselect),                                              //                                                     .chipselect
		.DIST2_s1_address                                                 (mm_interconnect_0_dist2_s1_address),                                                 //                                             DIST2_s1.address
		.DIST2_s1_write                                                   (mm_interconnect_0_dist2_s1_write),                                                   //                                                     .write
		.DIST2_s1_read                                                    (mm_interconnect_0_dist2_s1_read),                                                    //                                                     .read
		.DIST2_s1_readdata                                                (mm_interconnect_0_dist2_s1_readdata),                                                //                                                     .readdata
		.DIST2_s1_writedata                                               (mm_interconnect_0_dist2_s1_writedata),                                               //                                                     .writedata
		.DIST2_s1_begintransfer                                           (mm_interconnect_0_dist2_s1_begintransfer),                                           //                                                     .begintransfer
		.DIST2_s1_chipselect                                              (mm_interconnect_0_dist2_s1_chipselect),                                              //                                                     .chipselect
		.DIST3_s1_address                                                 (mm_interconnect_0_dist3_s1_address),                                                 //                                             DIST3_s1.address
		.DIST3_s1_write                                                   (mm_interconnect_0_dist3_s1_write),                                                   //                                                     .write
		.DIST3_s1_read                                                    (mm_interconnect_0_dist3_s1_read),                                                    //                                                     .read
		.DIST3_s1_readdata                                                (mm_interconnect_0_dist3_s1_readdata),                                                //                                                     .readdata
		.DIST3_s1_writedata                                               (mm_interconnect_0_dist3_s1_writedata),                                               //                                                     .writedata
		.DIST3_s1_begintransfer                                           (mm_interconnect_0_dist3_s1_begintransfer),                                           //                                                     .begintransfer
		.DIST3_s1_chipselect                                              (mm_interconnect_0_dist3_s1_chipselect),                                              //                                                     .chipselect
		.DIST4_s1_address                                                 (mm_interconnect_0_dist4_s1_address),                                                 //                                             DIST4_s1.address
		.DIST4_s1_write                                                   (mm_interconnect_0_dist4_s1_write),                                                   //                                                     .write
		.DIST4_s1_read                                                    (mm_interconnect_0_dist4_s1_read),                                                    //                                                     .read
		.DIST4_s1_readdata                                                (mm_interconnect_0_dist4_s1_readdata),                                                //                                                     .readdata
		.DIST4_s1_writedata                                               (mm_interconnect_0_dist4_s1_writedata),                                               //                                                     .writedata
		.DIST4_s1_begintransfer                                           (mm_interconnect_0_dist4_s1_begintransfer),                                           //                                                     .begintransfer
		.DIST4_s1_chipselect                                              (mm_interconnect_0_dist4_s1_chipselect),                                              //                                                     .chipselect
		.DIST5_s1_address                                                 (mm_interconnect_0_dist5_s1_address),                                                 //                                             DIST5_s1.address
		.DIST5_s1_write                                                   (mm_interconnect_0_dist5_s1_write),                                                   //                                                     .write
		.DIST5_s1_read                                                    (mm_interconnect_0_dist5_s1_read),                                                    //                                                     .read
		.DIST5_s1_readdata                                                (mm_interconnect_0_dist5_s1_readdata),                                                //                                                     .readdata
		.DIST5_s1_writedata                                               (mm_interconnect_0_dist5_s1_writedata),                                               //                                                     .writedata
		.DIST5_s1_begintransfer                                           (mm_interconnect_0_dist5_s1_begintransfer),                                           //                                                     .begintransfer
		.DIST5_s1_chipselect                                              (mm_interconnect_0_dist5_s1_chipselect),                                              //                                                     .chipselect
		.DIST6_s1_address                                                 (mm_interconnect_0_dist6_s1_address),                                                 //                                             DIST6_s1.address
		.DIST6_s1_write                                                   (mm_interconnect_0_dist6_s1_write),                                                   //                                                     .write
		.DIST6_s1_read                                                    (mm_interconnect_0_dist6_s1_read),                                                    //                                                     .read
		.DIST6_s1_readdata                                                (mm_interconnect_0_dist6_s1_readdata),                                                //                                                     .readdata
		.DIST6_s1_writedata                                               (mm_interconnect_0_dist6_s1_writedata),                                               //                                                     .writedata
		.DIST6_s1_begintransfer                                           (mm_interconnect_0_dist6_s1_begintransfer),                                           //                                                     .begintransfer
		.DIST6_s1_chipselect                                              (mm_interconnect_0_dist6_s1_chipselect),                                              //                                                     .chipselect
		.DIST7_s1_address                                                 (mm_interconnect_0_dist7_s1_address),                                                 //                                             DIST7_s1.address
		.DIST7_s1_write                                                   (mm_interconnect_0_dist7_s1_write),                                                   //                                                     .write
		.DIST7_s1_read                                                    (mm_interconnect_0_dist7_s1_read),                                                    //                                                     .read
		.DIST7_s1_readdata                                                (mm_interconnect_0_dist7_s1_readdata),                                                //                                                     .readdata
		.DIST7_s1_writedata                                               (mm_interconnect_0_dist7_s1_writedata),                                               //                                                     .writedata
		.DIST7_s1_begintransfer                                           (mm_interconnect_0_dist7_s1_begintransfer),                                           //                                                     .begintransfer
		.DIST7_s1_chipselect                                              (mm_interconnect_0_dist7_s1_chipselect),                                              //                                                     .chipselect
		.DIST8_s1_address                                                 (mm_interconnect_0_dist8_s1_address),                                                 //                                             DIST8_s1.address
		.DIST8_s1_write                                                   (mm_interconnect_0_dist8_s1_write),                                                   //                                                     .write
		.DIST8_s1_read                                                    (mm_interconnect_0_dist8_s1_read),                                                    //                                                     .read
		.DIST8_s1_readdata                                                (mm_interconnect_0_dist8_s1_readdata),                                                //                                                     .readdata
		.DIST8_s1_writedata                                               (mm_interconnect_0_dist8_s1_writedata),                                               //                                                     .writedata
		.DIST8_s1_begintransfer                                           (mm_interconnect_0_dist8_s1_begintransfer),                                           //                                                     .begintransfer
		.DIST8_s1_chipselect                                              (mm_interconnect_0_dist8_s1_chipselect),                                              //                                                     .chipselect
		.ENCODER_INT_s1_address                                           (mm_interconnect_0_encoder_int_s1_address),                                           //                                       ENCODER_INT_s1.address
		.ENCODER_INT_s1_write                                             (mm_interconnect_0_encoder_int_s1_write),                                             //                                                     .write
		.ENCODER_INT_s1_readdata                                          (mm_interconnect_0_encoder_int_s1_readdata),                                          //                                                     .readdata
		.ENCODER_INT_s1_writedata                                         (mm_interconnect_0_encoder_int_s1_writedata),                                         //                                                     .writedata
		.ENCODER_INT_s1_chipselect                                        (mm_interconnect_0_encoder_int_s1_chipselect),                                        //                                                     .chipselect
		.ENCODER_NORMAL_s1_address                                        (mm_interconnect_0_encoder_normal_s1_address),                                        //                                    ENCODER_NORMAL_s1.address
		.ENCODER_NORMAL_s1_readdata                                       (mm_interconnect_0_encoder_normal_s1_readdata),                                       //                                                     .readdata
		.EPCS_epcs_control_port_address                                   (mm_interconnect_0_epcs_epcs_control_port_address),                                   //                               EPCS_epcs_control_port.address
		.EPCS_epcs_control_port_write                                     (mm_interconnect_0_epcs_epcs_control_port_write),                                     //                                                     .write
		.EPCS_epcs_control_port_read                                      (mm_interconnect_0_epcs_epcs_control_port_read),                                      //                                                     .read
		.EPCS_epcs_control_port_readdata                                  (mm_interconnect_0_epcs_epcs_control_port_readdata),                                  //                                                     .readdata
		.EPCS_epcs_control_port_writedata                                 (mm_interconnect_0_epcs_epcs_control_port_writedata),                                 //                                                     .writedata
		.EPCS_epcs_control_port_chipselect                                (mm_interconnect_0_epcs_epcs_control_port_chipselect),                                //                                                     .chipselect
		.FLAG_I2C_s1_address                                              (mm_interconnect_0_flag_i2c_s1_address),                                              //                                          FLAG_I2C_s1.address
		.FLAG_I2C_s1_readdata                                             (mm_interconnect_0_flag_i2c_s1_readdata),                                             //                                                     .readdata
		.GPS_s1_address                                                   (mm_interconnect_0_gps_s1_address),                                                   //                                               GPS_s1.address
		.GPS_s1_write                                                     (mm_interconnect_0_gps_s1_write),                                                     //                                                     .write
		.GPS_s1_read                                                      (mm_interconnect_0_gps_s1_read),                                                      //                                                     .read
		.GPS_s1_readdata                                                  (mm_interconnect_0_gps_s1_readdata),                                                  //                                                     .readdata
		.GPS_s1_writedata                                                 (mm_interconnect_0_gps_s1_writedata),                                                 //                                                     .writedata
		.GPS_s1_begintransfer                                             (mm_interconnect_0_gps_s1_begintransfer),                                             //                                                     .begintransfer
		.GPS_s1_chipselect                                                (mm_interconnect_0_gps_s1_chipselect),                                                //                                                     .chipselect
		.JTAG_avalon_jtag_slave_address                                   (mm_interconnect_0_jtag_avalon_jtag_slave_address),                                   //                               JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write                                     (mm_interconnect_0_jtag_avalon_jtag_slave_write),                                     //                                                     .write
		.JTAG_avalon_jtag_slave_read                                      (mm_interconnect_0_jtag_avalon_jtag_slave_read),                                      //                                                     .read
		.JTAG_avalon_jtag_slave_readdata                                  (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),                                  //                                                     .readdata
		.JTAG_avalon_jtag_slave_writedata                                 (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),                                 //                                                     .writedata
		.JTAG_avalon_jtag_slave_waitrequest                               (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest),                               //                                                     .waitrequest
		.JTAG_avalon_jtag_slave_chipselect                                (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),                                //                                                     .chipselect
		.KEY_s1_address                                                   (mm_interconnect_0_key_s1_address),                                                   //                                               KEY_s1.address
		.KEY_s1_write                                                     (mm_interconnect_0_key_s1_write),                                                     //                                                     .write
		.KEY_s1_readdata                                                  (mm_interconnect_0_key_s1_readdata),                                                  //                                                     .readdata
		.KEY_s1_writedata                                                 (mm_interconnect_0_key_s1_writedata),                                                 //                                                     .writedata
		.KEY_s1_chipselect                                                (mm_interconnect_0_key_s1_chipselect),                                                //                                                     .chipselect
		.LED_s1_address                                                   (mm_interconnect_0_led_s1_address),                                                   //                                               LED_s1.address
		.LED_s1_write                                                     (mm_interconnect_0_led_s1_write),                                                     //                                                     .write
		.LED_s1_readdata                                                  (mm_interconnect_0_led_s1_readdata),                                                  //                                                     .readdata
		.LED_s1_writedata                                                 (mm_interconnect_0_led_s1_writedata),                                                 //                                                     .writedata
		.LED_s1_chipselect                                                (mm_interconnect_0_led_s1_chipselect),                                                //                                                     .chipselect
		.MOTORES_s1_address                                               (mm_interconnect_0_motores_s1_address),                                               //                                           MOTORES_s1.address
		.MOTORES_s1_write                                                 (mm_interconnect_0_motores_s1_write),                                                 //                                                     .write
		.MOTORES_s1_readdata                                              (mm_interconnect_0_motores_s1_readdata),                                              //                                                     .readdata
		.MOTORES_s1_writedata                                             (mm_interconnect_0_motores_s1_writedata),                                             //                                                     .writedata
		.MOTORES_s1_chipselect                                            (mm_interconnect_0_motores_s1_chipselect),                                            //                                                     .chipselect
		.PWM1_s1_address                                                  (mm_interconnect_0_pwm1_s1_address),                                                  //                                              PWM1_s1.address
		.PWM1_s1_write                                                    (mm_interconnect_0_pwm1_s1_write),                                                    //                                                     .write
		.PWM1_s1_readdata                                                 (mm_interconnect_0_pwm1_s1_readdata),                                                 //                                                     .readdata
		.PWM1_s1_writedata                                                (mm_interconnect_0_pwm1_s1_writedata),                                                //                                                     .writedata
		.PWM1_s1_chipselect                                               (mm_interconnect_0_pwm1_s1_chipselect),                                               //                                                     .chipselect
		.PWM2_s1_address                                                  (mm_interconnect_0_pwm2_s1_address),                                                  //                                              PWM2_s1.address
		.PWM2_s1_write                                                    (mm_interconnect_0_pwm2_s1_write),                                                    //                                                     .write
		.PWM2_s1_readdata                                                 (mm_interconnect_0_pwm2_s1_readdata),                                                 //                                                     .readdata
		.PWM2_s1_writedata                                                (mm_interconnect_0_pwm2_s1_writedata),                                                //                                                     .writedata
		.PWM2_s1_chipselect                                               (mm_interconnect_0_pwm2_s1_chipselect),                                               //                                                     .chipselect
		.SDRAM_s1_address                                                 (mm_interconnect_0_sdram_s1_address),                                                 //                                             SDRAM_s1.address
		.SDRAM_s1_write                                                   (mm_interconnect_0_sdram_s1_write),                                                   //                                                     .write
		.SDRAM_s1_read                                                    (mm_interconnect_0_sdram_s1_read),                                                    //                                                     .read
		.SDRAM_s1_readdata                                                (mm_interconnect_0_sdram_s1_readdata),                                                //                                                     .readdata
		.SDRAM_s1_writedata                                               (mm_interconnect_0_sdram_s1_writedata),                                               //                                                     .writedata
		.SDRAM_s1_byteenable                                              (mm_interconnect_0_sdram_s1_byteenable),                                              //                                                     .byteenable
		.SDRAM_s1_readdatavalid                                           (mm_interconnect_0_sdram_s1_readdatavalid),                                           //                                                     .readdatavalid
		.SDRAM_s1_waitrequest                                             (mm_interconnect_0_sdram_s1_waitrequest),                                             //                                                     .waitrequest
		.SDRAM_s1_chipselect                                              (mm_interconnect_0_sdram_s1_chipselect),                                              //                                                     .chipselect
		.SW_s1_address                                                    (mm_interconnect_0_sw_s1_address),                                                    //                                                SW_s1.address
		.SW_s1_readdata                                                   (mm_interconnect_0_sw_s1_readdata),                                                   //                                                     .readdata
		.sys_id_control_slave_address                                     (mm_interconnect_0_sys_id_control_slave_address),                                     //                                 sys_id_control_slave.address
		.sys_id_control_slave_readdata                                    (mm_interconnect_0_sys_id_control_slave_readdata),                                    //                                                     .readdata
		.sys_pll_pll_slave_address                                        (mm_interconnect_0_sys_pll_pll_slave_address),                                        //                                    sys_pll_pll_slave.address
		.sys_pll_pll_slave_write                                          (mm_interconnect_0_sys_pll_pll_slave_write),                                          //                                                     .write
		.sys_pll_pll_slave_read                                           (mm_interconnect_0_sys_pll_pll_slave_read),                                           //                                                     .read
		.sys_pll_pll_slave_readdata                                       (mm_interconnect_0_sys_pll_pll_slave_readdata),                                       //                                                     .readdata
		.sys_pll_pll_slave_writedata                                      (mm_interconnect_0_sys_pll_pll_slave_writedata),                                      //                                                     .writedata
		.sys_timer_s1_address                                             (mm_interconnect_0_sys_timer_s1_address),                                             //                                         sys_timer_s1.address
		.sys_timer_s1_write                                               (mm_interconnect_0_sys_timer_s1_write),                                               //                                                     .write
		.sys_timer_s1_readdata                                            (mm_interconnect_0_sys_timer_s1_readdata),                                            //                                                     .readdata
		.sys_timer_s1_writedata                                           (mm_interconnect_0_sys_timer_s1_writedata),                                           //                                                     .writedata
		.sys_timer_s1_chipselect                                          (mm_interconnect_0_sys_timer_s1_chipselect),                                          //                                                     .chipselect
		.XBEE_s1_address                                                  (mm_interconnect_0_xbee_s1_address),                                                  //                                              XBEE_s1.address
		.XBEE_s1_write                                                    (mm_interconnect_0_xbee_s1_write),                                                    //                                                     .write
		.XBEE_s1_read                                                     (mm_interconnect_0_xbee_s1_read),                                                     //                                                     .read
		.XBEE_s1_readdata                                                 (mm_interconnect_0_xbee_s1_readdata),                                                 //                                                     .readdata
		.XBEE_s1_writedata                                                (mm_interconnect_0_xbee_s1_writedata),                                                //                                                     .writedata
		.XBEE_s1_begintransfer                                            (mm_interconnect_0_xbee_s1_begintransfer),                                            //                                                     .begintransfer
		.XBEE_s1_chipselect                                               (mm_interconnect_0_xbee_s1_chipselect)                                                //                                                     .chipselect
	);

	NIOS_irq_mapper irq_mapper (
		.clk            (sys_pll_c0_clk),                 //        clk.clk
		.reset          (rst_controller_reset_out_reset), //  clk_reset.reset
		.receiver0_irq  (irq_mapper_receiver0_irq),       //  receiver0.irq
		.receiver1_irq  (irq_mapper_receiver1_irq),       //  receiver1.irq
		.receiver2_irq  (irq_mapper_receiver2_irq),       //  receiver2.irq
		.receiver3_irq  (irq_mapper_receiver3_irq),       //  receiver3.irq
		.receiver4_irq  (irq_mapper_receiver4_irq),       //  receiver4.irq
		.receiver5_irq  (irq_mapper_receiver5_irq),       //  receiver5.irq
		.receiver6_irq  (irq_mapper_receiver6_irq),       //  receiver6.irq
		.receiver7_irq  (irq_mapper_receiver7_irq),       //  receiver7.irq
		.receiver8_irq  (irq_mapper_receiver8_irq),       //  receiver8.irq
		.receiver9_irq  (irq_mapper_receiver9_irq),       //  receiver9.irq
		.receiver10_irq (irq_mapper_receiver10_irq),      // receiver10.irq
		.receiver11_irq (irq_mapper_receiver11_irq),      // receiver11.irq
		.receiver12_irq (irq_mapper_receiver12_irq),      // receiver12.irq
		.receiver13_irq (irq_mapper_receiver13_irq),      // receiver13.irq
		.receiver14_irq (irq_mapper_receiver14_irq),      // receiver14.irq
		.receiver15_irq (irq_mapper_receiver15_irq),      // receiver15.irq
		.sender_irq     (cpu_d_irq_irq)                   //     sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.reset_in2      (rst_controller_002_reset_out_reset), // reset_in2.reset
		.reset_in3      (rst_controller_003_reset_out_reset), // reset_in3.reset
		.clk            (sys_pll_c0_clk),                     //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (4),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.reset_in2      (rst_controller_002_reset_out_reset), // reset_in2.reset
		.reset_in3      (rst_controller_003_reset_out_reset), // reset_in3.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
